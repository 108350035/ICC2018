module CHIP(clk, 
		reset, 
		cmd, 
		cmd_valid, 
             IROM_rd, 
		 IROM_A, 
		IROM_Q, 
             IRAM_valid, 
		IRAM_D, IRAM_A,
		     busy, done);
input clk;
input reset;
input [3:0] cmd;
input cmd_valid;
input [7:0] IROM_Q;
output IROM_rd;
output [5:0] IROM_A;
output IRAM_valid;
output [7:0] IRAM_D;
output [5:0] IRAM_A;
output busy;
output done;


wire C_clk;
wire C_reset;
wire [3:0] C_cmd;
wire C_cmd_valid;
wire [7:0] C_IROM_Q;
wire  C_IROM_rd;
wire [5:0] C_IROM_A;
wire  C_IRAM_valid;
wire [7:0] C_IRAM_D;
wire [5:0] C_IRAM_A;
wire  C_busy;
wire C_done;




wire BUF_clk;
CLKBUFX20 buf0(.A(C_clk),.Y(BUF_clk));

LCD_CTRL LCD_CTRL(.clk(BUF_clk), .reset(C_reset), 
		     .cmd(C_cmd), .cmd_valid(C_cmd_valid), 
                     .IROM_rd(C_IROM_rd), .IROM_A(C_IROM_A), .IROM_Q(C_IROM_Q), 
                     .IRAM_valid(C_IRAM_valid), .IRAM_D(C_IRAM_D), .IRAM_A(C_IRAM_A),
		     .busy(C_busy), .done(C_done));


// Input Pads
PDUSDGZ I_CLK(.PAD(clk), .C(C_clk));
PDUSDGZ I_RESET(.PAD(reset), .C(C_reset));
PDUSDGZ I_CMD_V  (.PAD(cmd_valid),  .C(C_cmd_valid));
PDUSDGZ I_CMD_0  (.PAD(cmd[0]),  .C(C_cmd[0]));
PDUSDGZ I_CMD_1  (.PAD(cmd[1]),  .C(C_cmd[1]));
PDUSDGZ I_CMD_2  (.PAD(cmd[2]),  .C(C_cmd[2]));
PDUSDGZ I_CMD_3  (.PAD(cmd[3]),  .C(C_cmd[3]));
PDUSDGZ I_ROMQ0  (.PAD(IROM_Q[0]),  .C(C_IROM_Q[0]));
PDUSDGZ I_ROMQ1  (.PAD(IROM_Q[1]),  .C(C_IROM_Q[1]));
PDUSDGZ I_ROMQ2  (.PAD(IROM_Q[2]),  .C(C_IROM_Q[2]));
PDUSDGZ I_ROMQ3  (.PAD(IROM_Q[3]),  .C(C_IROM_Q[3]));
PDUSDGZ I_ROMQ4  (.PAD(IROM_Q[4]),  .C(C_IROM_Q[4]));
PDUSDGZ I_ROMQ5  (.PAD(IROM_Q[5]),  .C(C_IROM_Q[5]));
PDUSDGZ I_ROMQ6  (.PAD(IROM_Q[6]),  .C(C_IROM_Q[6]));
PDUSDGZ I_ROMQ7  (.PAD(IROM_Q[7]),  .C(C_IROM_Q[7]));


// Output Pads
PDD08SDGZ O_BUSY  (.OEN(1'b0), .I(C_busy),  .PAD(busy),  .C());
PDD08SDGZ O_DONE  (.OEN(1'b0), .I(C_done),  .PAD(done),  .C());
PDD08SDGZ O_IRAM_V  (.OEN(1'b0), .I(C_IRAM_valid),  .PAD(IRAM_valid),  .C());
PDD08SDGZ O_IRAMD0  (.OEN(1'b0), .I(C_IRAM_D[0]),  .PAD(IRAM_D[0]),  .C());
PDD08SDGZ O_IRAMD1  (.OEN(1'b0), .I(C_IRAM_D[1]),  .PAD(IRAM_D[1]),  .C());
PDD08SDGZ O_IRAMD2  (.OEN(1'b0), .I(C_IRAM_D[2]),  .PAD(IRAM_D[2]),  .C());
PDD08SDGZ O_IRAMD3  (.OEN(1'b0), .I(C_IRAM_D[3]),  .PAD(IRAM_D[3]),  .C());
PDD08SDGZ O_IRAMD4  (.OEN(1'b0), .I(C_IRAM_D[4]),  .PAD(IRAM_D[4]),  .C());
PDD08SDGZ O_IRAMD5  (.OEN(1'b0), .I(C_IRAM_D[5]),  .PAD(IRAM_D[5]),  .C());
PDD08SDGZ O_IRAMD6  (.OEN(1'b0), .I(C_IRAM_D[6]),  .PAD(IRAM_D[6]),  .C());
PDD08SDGZ O_IRAMD7  (.OEN(1'b0), .I(C_IRAM_D[7]),  .PAD(IRAM_D[7]),  .C());
PDD08SDGZ O_IRAMA0  (.OEN(1'b0), .I(C_IRAM_A[0]),  .PAD(IRAM_A[0]),  .C());
PDD08SDGZ O_IRAMA1  (.OEN(1'b0), .I(C_IRAM_A[1]),  .PAD(IRAM_A[1]),  .C());
PDD08SDGZ O_IRAMA2  (.OEN(1'b0), .I(C_IRAM_A[2]),  .PAD(IRAM_A[2]),  .C());
PDD08SDGZ O_IRAMA3  (.OEN(1'b0), .I(C_IRAM_A[3]),  .PAD(IRAM_A[3]),  .C());
PDD08SDGZ O_IRAMA4  (.OEN(1'b0), .I(C_IRAM_A[4]),  .PAD(IRAM_A[4]),  .C());
PDD08SDGZ O_IRAMA5  (.OEN(1'b0), .I(C_IRAM_A[5]),  .PAD(IRAM_A[5]),  .C());
PDD08SDGZ O_IROMA0  (.OEN(1'b0), .I(C_IROM_A[0]),  .PAD(IROM_A[0]),  .C());
PDD08SDGZ O_IROMA1  (.OEN(1'b0), .I(C_IROM_A[1]),  .PAD(IROM_A[1]),  .C());
PDD08SDGZ O_IROMA2  (.OEN(1'b0), .I(C_IROM_A[2]),  .PAD(IROM_A[2]),  .C());
PDD08SDGZ O_IROMA3  (.OEN(1'b0), .I(C_IROM_A[3]),  .PAD(IROM_A[3]),  .C());
PDD08SDGZ O_IROMA4  (.OEN(1'b0), .I(C_IROM_A[4]),  .PAD(IROM_A[4]),  .C());
PDD08SDGZ O_IROMA5  (.OEN(1'b0), .I(C_IROM_A[5]),  .PAD(IROM_A[5]),  .C());
PDD08SDGZ O_IROMRD  (.OEN(1'b0), .I(C_IROM_rd),  .PAD(IROM_rd),  .C());
// IO power 
PVDD2DGZ VDDP0 ();
PVSS2DGZ GNDP0 ();
PVDD2DGZ VDDP1 ();
PVSS2DGZ GNDP1 ();
PVDD2DGZ VDDP2 ();
PVSS2DGZ GNDP2 ();
PVDD2DGZ VDDP3 ();
PVSS2DGZ GNDP3 ();



// Core power
PVDD1DGZ VDDC0 ();
PVSS1DGZ GNDC0 ();
PVDD1DGZ VDDC1 ();
PVSS1DGZ GNDC1 ();
PVDD1DGZ VDDC2 ();
PVSS1DGZ GNDC2 ();
PVDD1DGZ VDDC3 ();
PVSS1DGZ GNDC3 ();



endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : O-2018.06-SP1
// Date      : Thu Dec 11 09:54:28 2025
/////////////////////////////////////////////////////////////


module LCD_CTRL ( clk, reset, cmd, cmd_valid, IROM_Q, IROM_rd, IROM_A, 
        IRAM_valid, IRAM_D, IRAM_A, busy, done );
  input [3:0] cmd;
  input [7:0] IROM_Q;
  output [5:0] IROM_A;
  output [7:0] IRAM_D;
  output [5:0] IRAM_A;
  input clk, reset, cmd_valid;
  output IROM_rd, IRAM_valid, busy, done;
  wire   in_valid, in_done, N2755, N2756, N2757, N2758, N2759, N2760, N2763,
         N2765, N2766, N2771, N2772, N2773, N2774, N2775, N2776, N2779, N2780,
         N2781, N2782, N2783, N2784, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         DP_OP_2677J1_122_9848_n30, DP_OP_2677J1_122_9848_n27,
         DP_OP_2677J1_122_9848_n26, DP_OP_2677J1_122_9848_n25,
         DP_OP_2677J1_122_9848_n24, DP_OP_2677J1_122_9848_n23,
         DP_OP_2677J1_122_9848_n22, DP_OP_2677J1_122_9848_n21,
         DP_OP_2677J1_122_9848_n20, DP_OP_2677J1_122_9848_n19,
         DP_OP_2677J1_122_9848_n18, DP_OP_2677J1_122_9848_n17,
         DP_OP_2677J1_122_9848_n16, DP_OP_2677J1_122_9848_n15,
         DP_OP_2677J1_122_9848_n14, DP_OP_2677J1_122_9848_n13,
         DP_OP_2677J1_122_9848_n12, DP_OP_2677J1_122_9848_n11,
         DP_OP_2677J1_122_9848_n10, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602;
  wire   [5:3] op4;
  wire   [2:0] op2;
  wire   [511:0] image_data;
  wire   [1:0] cs;
  wire   [3:0] cmd_reg;

  DFFSX1 cmd_reg_reg_3_ ( .D(n3337), .CK(clk), .SN(n8583), .QN(cmd_reg[3]) );
  DFFSX1 cmd_reg_reg_2_ ( .D(n3336), .CK(clk), .SN(n8578), .Q(n8532), .QN(
        cmd_reg[2]) );
  DFFSX1 cmd_reg_reg_1_ ( .D(n3335), .CK(clk), .SN(n8571), .QN(cmd_reg[1]) );
  DFFSX1 cmd_reg_reg_0_ ( .D(n3334), .CK(clk), .SN(n8595), .Q(n8531), .QN(
        cmd_reg[0]) );
  DFFSX1 in_done_reg ( .D(n3329), .CK(clk), .SN(n8590), .QN(in_done) );
  DFFSX1 y_cal_reg_1_ ( .D(n3325), .CK(clk), .SN(n8594), .Q(n8518), .QN(op4[4]) );
  DFFSX1 x_cal_reg_1_ ( .D(n3323), .CK(clk), .SN(n8586), .Q(n8530), .QN(op2[1]) );
  DFFSX1 in_valid_reg ( .D(n8566), .CK(clk), .SN(n8592), .Q(n8523), .QN(
        in_valid) );
  DFFSX1 image_data_reg_63__7_ ( .D(n3319), .CK(clk), .SN(n8573), .QN(
        image_data[511]) );
  DFFSX1 image_data_reg_63__6_ ( .D(n3318), .CK(clk), .SN(n8598), .QN(
        image_data[510]) );
  DFFSX1 image_data_reg_63__5_ ( .D(n3317), .CK(clk), .SN(n8601), .QN(
        image_data[509]) );
  DFFSX1 image_data_reg_63__4_ ( .D(n3316), .CK(clk), .SN(n8597), .QN(
        image_data[508]) );
  DFFSX1 image_data_reg_63__3_ ( .D(n3315), .CK(clk), .SN(n8585), .QN(
        image_data[507]) );
  DFFSX1 image_data_reg_63__2_ ( .D(n3314), .CK(clk), .SN(n8584), .QN(
        image_data[506]) );
  DFFSX1 image_data_reg_63__1_ ( .D(n3313), .CK(clk), .SN(n8583), .QN(
        image_data[505]) );
  DFFSX1 image_data_reg_63__0_ ( .D(n3312), .CK(clk), .SN(n8576), .QN(
        image_data[504]) );
  DFFSX1 image_data_reg_62__7_ ( .D(n3311), .CK(clk), .SN(n8577), .QN(
        image_data[503]) );
  DFFSX1 image_data_reg_62__6_ ( .D(n3310), .CK(clk), .SN(n8578), .QN(
        image_data[502]) );
  DFFSX1 image_data_reg_62__5_ ( .D(n3309), .CK(clk), .SN(n8579), .QN(
        image_data[501]) );
  DFFSX1 image_data_reg_62__4_ ( .D(n3308), .CK(clk), .SN(n8580), .QN(
        image_data[500]) );
  DFFSX1 image_data_reg_62__3_ ( .D(n3307), .CK(clk), .SN(n8583), .QN(
        image_data[499]) );
  DFFSX1 image_data_reg_62__2_ ( .D(n3306), .CK(clk), .SN(n8576), .QN(
        image_data[498]) );
  DFFSX1 image_data_reg_62__1_ ( .D(n3305), .CK(clk), .SN(n8577), .QN(
        image_data[497]) );
  DFFSX1 image_data_reg_62__0_ ( .D(n3304), .CK(clk), .SN(n8578), .QN(
        image_data[496]) );
  DFFSX1 image_data_reg_61__7_ ( .D(n3303), .CK(clk), .SN(n8579), .QN(
        image_data[495]) );
  DFFSX1 image_data_reg_61__6_ ( .D(n3302), .CK(clk), .SN(n8580), .QN(
        image_data[494]) );
  DFFSX1 image_data_reg_61__5_ ( .D(n3301), .CK(clk), .SN(n8594), .QN(
        image_data[493]) );
  DFFSX1 image_data_reg_61__4_ ( .D(n3300), .CK(clk), .SN(n8595), .QN(
        image_data[492]) );
  DFFSX1 image_data_reg_61__3_ ( .D(n3299), .CK(clk), .SN(n8586), .QN(
        image_data[491]) );
  DFFSX1 image_data_reg_61__2_ ( .D(n3298), .CK(clk), .SN(n8581), .QN(
        image_data[490]) );
  DFFSX1 image_data_reg_61__1_ ( .D(n3297), .CK(clk), .SN(n8582), .QN(
        image_data[489]) );
  DFFSX1 image_data_reg_61__0_ ( .D(n3296), .CK(clk), .SN(n8589), .QN(
        image_data[488]) );
  DFFSX1 image_data_reg_60__7_ ( .D(n3295), .CK(clk), .SN(n8594), .QN(
        image_data[487]) );
  DFFSX1 image_data_reg_60__6_ ( .D(n3294), .CK(clk), .SN(n8595), .QN(
        image_data[486]) );
  DFFSX1 image_data_reg_60__5_ ( .D(n3293), .CK(clk), .SN(n8586), .QN(
        image_data[485]) );
  DFFSX1 image_data_reg_60__4_ ( .D(n3292), .CK(clk), .SN(n8581), .QN(
        image_data[484]) );
  DFFSX1 image_data_reg_60__3_ ( .D(n3291), .CK(clk), .SN(n8582), .QN(
        image_data[483]) );
  DFFSX1 image_data_reg_60__2_ ( .D(n3290), .CK(clk), .SN(n8589), .QN(
        image_data[482]) );
  DFFSX1 image_data_reg_60__1_ ( .D(n3289), .CK(clk), .SN(n8592), .QN(
        image_data[481]) );
  DFFSX1 image_data_reg_60__0_ ( .D(n3288), .CK(clk), .SN(n8591), .QN(
        image_data[480]) );
  DFFSX1 image_data_reg_59__7_ ( .D(n3287), .CK(clk), .SN(n8590), .QN(
        image_data[479]) );
  DFFSX1 image_data_reg_59__6_ ( .D(n3286), .CK(clk), .SN(n8588), .QN(
        image_data[478]) );
  DFFSX1 image_data_reg_59__5_ ( .D(n3285), .CK(clk), .SN(n8587), .QN(
        image_data[477]) );
  DFFSX1 image_data_reg_59__4_ ( .D(n3284), .CK(clk), .SN(n8593), .QN(
        image_data[476]) );
  DFFSX1 image_data_reg_59__3_ ( .D(n3283), .CK(clk), .SN(n8570), .QN(
        image_data[475]) );
  DFFSX1 image_data_reg_59__2_ ( .D(n3282), .CK(clk), .SN(n8602), .QN(
        image_data[474]) );
  DFFSX1 image_data_reg_59__1_ ( .D(n3281), .CK(clk), .SN(n8575), .QN(
        image_data[473]) );
  DFFSX1 image_data_reg_59__0_ ( .D(n3280), .CK(clk), .SN(n8599), .QN(
        image_data[472]) );
  DFFSX1 image_data_reg_58__7_ ( .D(n3279), .CK(clk), .SN(n8572), .QN(
        image_data[471]) );
  DFFSX1 image_data_reg_58__6_ ( .D(n3278), .CK(clk), .SN(n8600), .Q(n8553), 
        .QN(image_data[470]) );
  DFFSX1 image_data_reg_58__5_ ( .D(n3277), .CK(clk), .SN(n8573), .QN(
        image_data[469]) );
  DFFSX1 image_data_reg_58__4_ ( .D(n3276), .CK(clk), .SN(n8598), .QN(
        image_data[468]) );
  DFFSX1 image_data_reg_58__3_ ( .D(n3275), .CK(clk), .SN(n8601), .QN(
        image_data[467]) );
  DFFSX1 image_data_reg_58__2_ ( .D(n3274), .CK(clk), .SN(n8597), .Q(n8556), 
        .QN(image_data[466]) );
  DFFSX1 image_data_reg_58__1_ ( .D(n3273), .CK(clk), .SN(n8585), .QN(
        image_data[465]) );
  DFFSX1 image_data_reg_58__0_ ( .D(n3272), .CK(clk), .SN(n8584), .QN(
        image_data[464]) );
  DFFSX1 image_data_reg_57__7_ ( .D(n3271), .CK(clk), .SN(n8578), .QN(
        image_data[463]) );
  DFFSX1 image_data_reg_57__6_ ( .D(n3270), .CK(clk), .SN(n8579), .QN(
        image_data[462]) );
  DFFSX1 image_data_reg_57__5_ ( .D(n3269), .CK(clk), .SN(n8580), .QN(
        image_data[461]) );
  DFFSX1 image_data_reg_57__4_ ( .D(n3268), .CK(clk), .SN(n8594), .QN(
        image_data[460]) );
  DFFSX1 image_data_reg_57__3_ ( .D(n3267), .CK(clk), .SN(n8595), .QN(
        image_data[459]) );
  DFFSX1 image_data_reg_57__2_ ( .D(n3266), .CK(clk), .SN(n8586), .QN(
        image_data[458]) );
  DFFSX1 image_data_reg_57__1_ ( .D(n3265), .CK(clk), .SN(n8581), .QN(
        image_data[457]) );
  DFFSX1 image_data_reg_57__0_ ( .D(n3264), .CK(clk), .SN(n8582), .QN(
        image_data[456]) );
  DFFSX1 image_data_reg_56__7_ ( .D(n3263), .CK(clk), .SN(n8589), .QN(
        image_data[455]) );
  DFFSX1 image_data_reg_56__6_ ( .D(n3262), .CK(clk), .SN(n8592), .QN(
        image_data[454]) );
  DFFSX1 image_data_reg_56__5_ ( .D(n3261), .CK(clk), .SN(n8591), .QN(
        image_data[453]) );
  DFFSX1 image_data_reg_56__4_ ( .D(n3260), .CK(clk), .SN(n8590), .Q(n8557), 
        .QN(image_data[452]) );
  DFFSX1 image_data_reg_56__3_ ( .D(n3259), .CK(clk), .SN(n8570), .QN(
        image_data[451]) );
  DFFSX1 image_data_reg_56__2_ ( .D(n3258), .CK(clk), .SN(n8602), .QN(
        image_data[450]) );
  DFFSX1 image_data_reg_56__1_ ( .D(n3257), .CK(clk), .SN(n8575), .QN(
        image_data[449]) );
  DFFSX1 image_data_reg_56__0_ ( .D(n3256), .CK(clk), .SN(n8599), .QN(
        image_data[448]) );
  DFFSX1 image_data_reg_55__7_ ( .D(n3255), .CK(clk), .SN(n8572), .QN(
        image_data[447]) );
  DFFSX1 image_data_reg_55__6_ ( .D(n3254), .CK(clk), .SN(n8600), .QN(
        image_data[446]) );
  DFFSX1 image_data_reg_55__5_ ( .D(n3253), .CK(clk), .SN(n8573), .QN(
        image_data[445]) );
  DFFSX1 image_data_reg_55__4_ ( .D(n3252), .CK(clk), .SN(n8598), .QN(
        image_data[444]) );
  DFFSX1 image_data_reg_55__3_ ( .D(n3251), .CK(clk), .SN(n8601), .QN(
        image_data[443]) );
  DFFSX1 image_data_reg_55__2_ ( .D(n3250), .CK(clk), .SN(n8597), .QN(
        image_data[442]) );
  DFFSX1 image_data_reg_55__1_ ( .D(n3249), .CK(clk), .SN(n8585), .QN(
        image_data[441]) );
  DFFSX1 image_data_reg_55__0_ ( .D(n3248), .CK(clk), .SN(n8584), .QN(
        image_data[440]) );
  DFFSX1 image_data_reg_54__7_ ( .D(n3247), .CK(clk), .SN(n8581), .QN(
        image_data[439]) );
  DFFSX1 image_data_reg_54__6_ ( .D(n3246), .CK(clk), .SN(n8582), .QN(
        image_data[438]) );
  DFFSX1 image_data_reg_54__5_ ( .D(n3245), .CK(clk), .SN(n8589), .QN(
        image_data[437]) );
  DFFSX1 image_data_reg_54__4_ ( .D(n3244), .CK(clk), .SN(n8592), .QN(
        image_data[436]) );
  DFFSX1 image_data_reg_54__3_ ( .D(n3243), .CK(clk), .SN(n8591), .QN(
        image_data[435]) );
  DFFSX1 image_data_reg_54__2_ ( .D(n3242), .CK(clk), .SN(n8590), .QN(
        image_data[434]) );
  DFFSX1 image_data_reg_54__1_ ( .D(n3241), .CK(clk), .SN(n8588), .QN(
        image_data[433]) );
  DFFSX1 image_data_reg_54__0_ ( .D(n3240), .CK(clk), .SN(n8587), .QN(
        image_data[432]) );
  DFFSX1 image_data_reg_53__7_ ( .D(n3239), .CK(clk), .SN(n8593), .QN(
        image_data[431]) );
  DFFSX1 image_data_reg_53__6_ ( .D(n3238), .CK(clk), .SN(n8579), .QN(
        image_data[430]) );
  DFFSX1 image_data_reg_53__5_ ( .D(n3237), .CK(clk), .SN(n8595), .QN(
        image_data[429]) );
  DFFSX1 image_data_reg_53__4_ ( .D(n3236), .CK(clk), .SN(n8571), .QN(
        image_data[428]) );
  DFFSX1 image_data_reg_53__3_ ( .D(n3235), .CK(clk), .SN(n8587), .QN(
        image_data[427]) );
  DFFSX1 image_data_reg_53__2_ ( .D(n3234), .CK(clk), .SN(n8576), .QN(
        image_data[426]) );
  DFFSX1 image_data_reg_53__1_ ( .D(n3233), .CK(clk), .SN(n8598), .QN(
        image_data[425]) );
  DFFSX1 image_data_reg_53__0_ ( .D(n3232), .CK(clk), .SN(n8587), .QN(
        image_data[424]) );
  DFFSX1 image_data_reg_52__7_ ( .D(n3231), .CK(clk), .SN(n8576), .QN(
        image_data[423]) );
  DFFSX1 image_data_reg_52__6_ ( .D(n3230), .CK(clk), .SN(n8574), .QN(
        image_data[422]) );
  DFFSX1 image_data_reg_52__5_ ( .D(n3229), .CK(clk), .SN(n8570), .QN(
        image_data[421]) );
  DFFSX1 image_data_reg_52__4_ ( .D(n3228), .CK(clk), .SN(n8586), .QN(
        image_data[420]) );
  DFFSX1 image_data_reg_52__3_ ( .D(n3227), .CK(clk), .SN(n8584), .QN(
        image_data[419]) );
  DFFSX1 image_data_reg_52__2_ ( .D(n3226), .CK(clk), .SN(n8571), .QN(
        image_data[418]) );
  DFFSX1 image_data_reg_52__1_ ( .D(n3225), .CK(clk), .SN(n8580), .QN(
        image_data[417]) );
  DFFSX1 image_data_reg_52__0_ ( .D(n3224), .CK(clk), .SN(n8575), .QN(
        image_data[416]) );
  DFFSX1 image_data_reg_51__7_ ( .D(n3223), .CK(clk), .SN(n8573), .QN(
        image_data[415]) );
  DFFSX1 image_data_reg_51__6_ ( .D(n3222), .CK(clk), .SN(n8598), .QN(
        image_data[414]) );
  DFFSX1 image_data_reg_51__5_ ( .D(n3221), .CK(clk), .SN(n8601), .QN(
        image_data[413]) );
  DFFSX1 image_data_reg_51__4_ ( .D(n3220), .CK(clk), .SN(n8597), .QN(
        image_data[412]) );
  DFFSX1 image_data_reg_51__3_ ( .D(n3219), .CK(clk), .SN(n8585), .QN(
        image_data[411]) );
  DFFSX1 image_data_reg_51__2_ ( .D(n3218), .CK(clk), .SN(n8584), .Q(n8558), 
        .QN(image_data[410]) );
  DFFSX1 image_data_reg_51__1_ ( .D(n3217), .CK(clk), .SN(n8583), .QN(
        image_data[409]) );
  DFFSX1 image_data_reg_51__0_ ( .D(n3216), .CK(clk), .SN(n8576), .QN(
        image_data[408]) );
  DFFSX1 image_data_reg_50__7_ ( .D(n3215), .CK(clk), .SN(n8577), .QN(
        image_data[407]) );
  DFFSX1 image_data_reg_50__6_ ( .D(n3214), .CK(clk), .SN(n8578), .QN(
        image_data[406]) );
  DFFSX1 image_data_reg_50__5_ ( .D(n3213), .CK(clk), .SN(n8579), .QN(
        image_data[405]) );
  DFFSX1 image_data_reg_50__4_ ( .D(n3212), .CK(clk), .SN(n8580), .QN(
        image_data[404]) );
  DFFSX1 image_data_reg_50__3_ ( .D(n3211), .CK(clk), .SN(n8594), .QN(
        image_data[403]) );
  DFFSX1 image_data_reg_50__2_ ( .D(n3210), .CK(clk), .SN(n8595), .QN(
        image_data[402]) );
  DFFSX1 image_data_reg_50__1_ ( .D(n3209), .CK(clk), .SN(n8588), .QN(
        image_data[401]) );
  DFFSX1 image_data_reg_50__0_ ( .D(n3208), .CK(clk), .SN(n8588), .QN(
        image_data[400]) );
  DFFSX1 image_data_reg_49__7_ ( .D(n3207), .CK(clk), .SN(n8597), .QN(
        image_data[399]) );
  DFFSX1 image_data_reg_49__6_ ( .D(n3206), .CK(clk), .SN(n8579), .QN(
        image_data[398]) );
  DFFSX1 image_data_reg_49__5_ ( .D(n3205), .CK(clk), .SN(n8578), .QN(
        image_data[397]) );
  DFFSX1 image_data_reg_49__4_ ( .D(n3204), .CK(clk), .SN(n8570), .QN(
        image_data[396]) );
  DFFSX1 image_data_reg_49__3_ ( .D(n3203), .CK(clk), .SN(n8587), .QN(
        image_data[395]) );
  DFFSX1 image_data_reg_49__2_ ( .D(n3202), .CK(clk), .SN(n8583), .QN(
        image_data[394]) );
  DFFSX1 image_data_reg_49__1_ ( .D(n3201), .CK(clk), .SN(n8587), .QN(
        image_data[393]) );
  DFFSX1 image_data_reg_49__0_ ( .D(n3200), .CK(clk), .SN(n8578), .QN(
        image_data[392]) );
  DFFSX1 image_data_reg_48__7_ ( .D(n3199), .CK(clk), .SN(n8587), .QN(
        image_data[391]) );
  DFFSX1 image_data_reg_48__6_ ( .D(n3198), .CK(clk), .SN(n8593), .QN(
        image_data[390]) );
  DFFSX1 image_data_reg_48__5_ ( .D(n3197), .CK(clk), .SN(n8583), .QN(
        image_data[389]) );
  DFFSX1 image_data_reg_48__4_ ( .D(n3196), .CK(clk), .SN(n8578), .QN(
        image_data[388]) );
  DFFSX1 image_data_reg_48__3_ ( .D(n3195), .CK(clk), .SN(n8571), .QN(
        image_data[387]) );
  DFFSX1 image_data_reg_48__2_ ( .D(n3194), .CK(clk), .SN(n8595), .QN(
        image_data[386]) );
  DFFSX1 image_data_reg_48__1_ ( .D(n3193), .CK(clk), .SN(n8574), .QN(
        image_data[385]) );
  DFFSX1 image_data_reg_48__0_ ( .D(n3192), .CK(clk), .SN(n8596), .Q(n8559), 
        .QN(image_data[384]) );
  DFFSX1 image_data_reg_47__7_ ( .D(n3191), .CK(clk), .SN(n8570), .QN(
        image_data[383]) );
  DFFSX1 image_data_reg_47__6_ ( .D(n3190), .CK(clk), .SN(n8602), .QN(
        image_data[382]) );
  DFFSX1 image_data_reg_47__5_ ( .D(n3189), .CK(clk), .SN(n8575), .QN(
        image_data[381]) );
  DFFSX1 image_data_reg_47__4_ ( .D(n3188), .CK(clk), .SN(n8599), .QN(
        image_data[380]) );
  DFFSX1 image_data_reg_47__3_ ( .D(n3187), .CK(clk), .SN(n8572), .QN(
        image_data[379]) );
  DFFSX1 image_data_reg_47__2_ ( .D(n3186), .CK(clk), .SN(n8600), .QN(
        image_data[378]) );
  DFFSX1 image_data_reg_47__1_ ( .D(n3185), .CK(clk), .SN(n8573), .QN(
        image_data[377]) );
  DFFSX1 image_data_reg_47__0_ ( .D(n3184), .CK(clk), .SN(n8598), .QN(
        image_data[376]) );
  DFFSX1 image_data_reg_46__7_ ( .D(n3183), .CK(clk), .SN(n8601), .QN(
        image_data[375]) );
  DFFSX1 image_data_reg_46__6_ ( .D(n3182), .CK(clk), .SN(n8597), .QN(
        image_data[374]) );
  DFFSX1 image_data_reg_46__5_ ( .D(n3181), .CK(clk), .SN(n8585), .QN(
        image_data[373]) );
  DFFSX1 image_data_reg_46__4_ ( .D(n3180), .CK(clk), .SN(n8584), .QN(
        image_data[372]) );
  DFFSX1 image_data_reg_46__3_ ( .D(n3179), .CK(clk), .SN(n8583), .QN(
        image_data[371]) );
  DFFSX1 image_data_reg_46__2_ ( .D(n3178), .CK(clk), .SN(n8576), .Q(n8539), 
        .QN(image_data[370]) );
  DFFSX1 image_data_reg_46__1_ ( .D(n3177), .CK(clk), .SN(n8577), .QN(
        image_data[369]) );
  DFFSX1 image_data_reg_46__0_ ( .D(n3176), .CK(clk), .SN(n8578), .QN(
        image_data[368]) );
  DFFSX1 image_data_reg_45__7_ ( .D(n3175), .CK(clk), .SN(n8574), .QN(
        image_data[367]) );
  DFFSX1 image_data_reg_45__6_ ( .D(n3174), .CK(clk), .SN(n8578), .QN(
        image_data[366]) );
  DFFSX1 image_data_reg_45__5_ ( .D(n3173), .CK(clk), .SN(n8595), .QN(
        image_data[365]) );
  DFFSX1 image_data_reg_45__4_ ( .D(n3172), .CK(clk), .SN(n8576), .QN(
        image_data[364]) );
  DFFSX1 image_data_reg_45__3_ ( .D(n3171), .CK(clk), .SN(n8585), .Q(n8540), 
        .QN(image_data[363]) );
  DFFSX1 image_data_reg_45__2_ ( .D(n3170), .CK(clk), .SN(n8595), .QN(
        image_data[362]) );
  DFFSX1 image_data_reg_45__1_ ( .D(n3169), .CK(clk), .SN(n8579), .Q(n8541), 
        .QN(image_data[361]) );
  DFFSX1 image_data_reg_45__0_ ( .D(n3168), .CK(clk), .SN(n8602), .QN(
        image_data[360]) );
  DFFSX1 image_data_reg_44__7_ ( .D(n3167), .CK(clk), .SN(n8593), .QN(
        image_data[359]) );
  DFFSX1 image_data_reg_44__6_ ( .D(n3166), .CK(clk), .SN(n8577), .QN(
        image_data[358]) );
  DFFSX1 image_data_reg_44__5_ ( .D(n3165), .CK(clk), .SN(n8593), .Q(n8535), 
        .QN(image_data[357]) );
  DFFSX1 image_data_reg_44__4_ ( .D(n3164), .CK(clk), .SN(n8596), .QN(
        image_data[356]) );
  DFFSX1 image_data_reg_44__3_ ( .D(n3163), .CK(clk), .SN(n8588), .QN(
        image_data[355]) );
  DFFSX1 image_data_reg_44__2_ ( .D(n3162), .CK(clk), .SN(n8601), .QN(
        image_data[354]) );
  DFFSX1 image_data_reg_44__1_ ( .D(n3161), .CK(clk), .SN(n8593), .QN(
        image_data[353]) );
  DFFSX1 image_data_reg_44__0_ ( .D(n3160), .CK(clk), .SN(n8577), .QN(
        image_data[352]) );
  DFFSX1 image_data_reg_43__7_ ( .D(n3159), .CK(clk), .SN(n8596), .QN(
        image_data[351]) );
  DFFSX1 image_data_reg_43__6_ ( .D(n3158), .CK(clk), .SN(n8578), .QN(
        image_data[350]) );
  DFFSX1 image_data_reg_43__5_ ( .D(n3157), .CK(clk), .SN(n8585), .QN(
        image_data[349]) );
  DFFSX1 image_data_reg_43__4_ ( .D(n3156), .CK(clk), .SN(n8594), .QN(
        image_data[348]) );
  DFFSX1 image_data_reg_43__3_ ( .D(n3155), .CK(clk), .SN(n8599), .QN(
        image_data[347]) );
  DFFSX1 image_data_reg_43__2_ ( .D(n3154), .CK(clk), .SN(n8592), .Q(n8542), 
        .QN(image_data[346]) );
  DFFSX1 image_data_reg_43__1_ ( .D(n3153), .CK(clk), .SN(n8584), .QN(
        image_data[345]) );
  DFFSX1 image_data_reg_43__0_ ( .D(n3152), .CK(clk), .SN(n8597), .QN(
        image_data[344]) );
  DFFSX1 image_data_reg_42__7_ ( .D(n3151), .CK(clk), .SN(n8591), .QN(
        image_data[343]) );
  DFFSX1 image_data_reg_42__6_ ( .D(n3150), .CK(clk), .SN(n8590), .Q(n8543), 
        .QN(image_data[342]) );
  DFFSX1 image_data_reg_42__5_ ( .D(n3149), .CK(clk), .SN(n8588), .QN(
        image_data[341]) );
  DFFSX1 image_data_reg_42__4_ ( .D(n3148), .CK(clk), .SN(n8587), .QN(
        image_data[340]) );
  DFFSX1 image_data_reg_42__3_ ( .D(n3147), .CK(clk), .SN(n8593), .QN(
        image_data[339]) );
  DFFSX1 image_data_reg_42__2_ ( .D(n3146), .CK(clk), .SN(n8577), .QN(
        image_data[338]) );
  DFFSX1 image_data_reg_42__1_ ( .D(n3145), .CK(clk), .SN(n8583), .QN(
        image_data[337]) );
  DFFSX1 image_data_reg_42__0_ ( .D(n3144), .CK(clk), .SN(n8571), .Q(n8544), 
        .QN(image_data[336]) );
  DFFSX1 image_data_reg_41__7_ ( .D(n3143), .CK(clk), .SN(n8579), .QN(
        image_data[335]) );
  DFFSX1 image_data_reg_41__6_ ( .D(n3142), .CK(clk), .SN(n8574), .QN(
        image_data[334]) );
  DFFSX1 image_data_reg_41__5_ ( .D(n3141), .CK(clk), .SN(n8596), .QN(
        image_data[333]) );
  DFFSX1 image_data_reg_41__4_ ( .D(n3140), .CK(clk), .SN(n8570), .QN(
        image_data[332]) );
  DFFSX1 image_data_reg_41__3_ ( .D(n3139), .CK(clk), .SN(n8586), .QN(
        image_data[331]) );
  DFFSX1 image_data_reg_41__2_ ( .D(n3138), .CK(clk), .SN(n8600), .QN(
        image_data[330]) );
  DFFSX1 image_data_reg_41__1_ ( .D(n3137), .CK(clk), .SN(n8590), .QN(
        image_data[329]) );
  DFFSX1 image_data_reg_41__0_ ( .D(n3136), .CK(clk), .SN(n8584), .QN(
        image_data[328]) );
  DFFSX1 image_data_reg_40__7_ ( .D(n3135), .CK(clk), .SN(n8571), .QN(
        image_data[327]) );
  DFFSX1 image_data_reg_40__6_ ( .D(n3134), .CK(clk), .SN(n8580), .Q(n8545), 
        .QN(image_data[326]) );
  DFFSX1 image_data_reg_40__5_ ( .D(n3133), .CK(clk), .SN(n8575), .QN(
        image_data[325]) );
  DFFSX1 image_data_reg_40__4_ ( .D(n3132), .CK(clk), .SN(n8589), .QN(
        image_data[324]) );
  DFFSX1 image_data_reg_40__3_ ( .D(n3131), .CK(clk), .SN(n8601), .QN(
        image_data[323]) );
  DFFSX1 image_data_reg_40__2_ ( .D(n3130), .CK(clk), .SN(n8593), .QN(
        image_data[322]) );
  DFFSX1 image_data_reg_40__1_ ( .D(n3129), .CK(clk), .SN(n8577), .QN(
        image_data[321]) );
  DFFSX1 image_data_reg_40__0_ ( .D(n3128), .CK(clk), .SN(n8596), .QN(
        image_data[320]) );
  DFFSX1 image_data_reg_39__7_ ( .D(n3127), .CK(clk), .SN(n8595), .QN(
        image_data[319]) );
  DFFSX1 image_data_reg_39__6_ ( .D(n3126), .CK(clk), .SN(n8571), .QN(
        image_data[318]) );
  DFFSX1 image_data_reg_39__5_ ( .D(n3125), .CK(clk), .SN(n8571), .QN(
        image_data[317]) );
  DFFSX1 image_data_reg_39__4_ ( .D(n3124), .CK(clk), .SN(n8577), .QN(
        image_data[316]) );
  DFFSX1 image_data_reg_39__3_ ( .D(n3123), .CK(clk), .SN(n8574), .QN(
        image_data[315]) );
  DFFSX1 image_data_reg_39__2_ ( .D(n3122), .CK(clk), .SN(n8596), .QN(
        image_data[314]) );
  DFFSX1 image_data_reg_39__1_ ( .D(n3121), .CK(clk), .SN(n8570), .QN(
        image_data[313]) );
  DFFSX1 image_data_reg_39__0_ ( .D(n3120), .CK(clk), .SN(n8602), .QN(
        image_data[312]) );
  DFFSX1 image_data_reg_38__7_ ( .D(n3119), .CK(clk), .SN(n8575), .QN(
        image_data[311]) );
  DFFSX1 image_data_reg_38__6_ ( .D(n3118), .CK(clk), .SN(n8599), .QN(
        image_data[310]) );
  DFFSX1 image_data_reg_38__5_ ( .D(n3117), .CK(clk), .SN(n8572), .QN(
        image_data[309]) );
  DFFSX1 image_data_reg_38__4_ ( .D(n3116), .CK(clk), .SN(n8600), .Q(n8536), 
        .QN(image_data[308]) );
  DFFSX1 image_data_reg_38__3_ ( .D(n3115), .CK(clk), .SN(n8597), .QN(
        image_data[307]) );
  DFFSX1 image_data_reg_38__2_ ( .D(n3114), .CK(clk), .SN(n8585), .QN(
        image_data[306]) );
  DFFSX1 image_data_reg_38__1_ ( .D(n3113), .CK(clk), .SN(n8584), .QN(
        image_data[305]) );
  DFFSX1 image_data_reg_38__0_ ( .D(n3112), .CK(clk), .SN(n8583), .QN(
        image_data[304]) );
  DFFSX1 image_data_reg_37__7_ ( .D(n3111), .CK(clk), .SN(n8576), .QN(
        image_data[303]) );
  DFFSX1 image_data_reg_37__6_ ( .D(n3110), .CK(clk), .SN(n8577), .QN(
        image_data[302]) );
  DFFSX1 image_data_reg_37__5_ ( .D(n3109), .CK(clk), .SN(n8578), .QN(
        image_data[301]) );
  DFFSX1 image_data_reg_37__4_ ( .D(n3108), .CK(clk), .SN(n8579), .QN(
        image_data[300]) );
  DFFSX1 image_data_reg_37__3_ ( .D(n3107), .CK(clk), .SN(n8580), .QN(
        image_data[299]) );
  DFFSX1 image_data_reg_37__2_ ( .D(n3106), .CK(clk), .SN(n8594), .QN(
        image_data[298]) );
  DFFSX1 image_data_reg_37__1_ ( .D(n3105), .CK(clk), .SN(n8595), .QN(
        image_data[297]) );
  DFFSX1 image_data_reg_37__0_ ( .D(n3104), .CK(clk), .SN(n8586), .QN(
        image_data[296]) );
  DFFSX1 image_data_reg_36__7_ ( .D(n3103), .CK(clk), .SN(n8592), .QN(
        image_data[295]) );
  DFFSX1 image_data_reg_36__6_ ( .D(n3102), .CK(clk), .SN(n8591), .QN(
        image_data[294]) );
  DFFSX1 image_data_reg_36__5_ ( .D(n3101), .CK(clk), .SN(n8590), .QN(
        image_data[293]) );
  DFFSX1 image_data_reg_36__4_ ( .D(n3100), .CK(clk), .SN(n8588), .QN(
        image_data[292]) );
  DFFSX1 image_data_reg_36__3_ ( .D(n3099), .CK(clk), .SN(n8587), .QN(
        image_data[291]) );
  DFFSX1 image_data_reg_36__2_ ( .D(n3098), .CK(clk), .SN(n8593), .QN(
        image_data[290]) );
  DFFSX1 image_data_reg_36__1_ ( .D(n3097), .CK(clk), .SN(n8578), .QN(
        image_data[289]) );
  DFFSX1 image_data_reg_36__0_ ( .D(n3096), .CK(clk), .SN(n8577), .QN(
        image_data[288]) );
  DFFSX1 image_data_reg_35__7_ ( .D(n3095), .CK(clk), .SN(n8571), .QN(
        image_data[287]) );
  DFFSX1 image_data_reg_35__6_ ( .D(n3094), .CK(clk), .SN(n8576), .QN(
        image_data[286]) );
  DFFSX1 image_data_reg_35__5_ ( .D(n3093), .CK(clk), .SN(n8574), .QN(
        image_data[285]) );
  DFFSX1 image_data_reg_35__4_ ( .D(n3092), .CK(clk), .SN(n8596), .QN(
        image_data[284]) );
  DFFSX1 image_data_reg_35__3_ ( .D(n3091), .CK(clk), .SN(n8595), .Q(n8546), 
        .QN(image_data[283]) );
  DFFSX1 image_data_reg_35__2_ ( .D(n3090), .CK(clk), .SN(n8586), .QN(
        image_data[282]) );
  DFFSX1 image_data_reg_35__1_ ( .D(n3089), .CK(clk), .SN(n8581), .QN(
        image_data[281]) );
  DFFSX1 image_data_reg_35__0_ ( .D(n3088), .CK(clk), .SN(n8582), .QN(
        image_data[280]) );
  DFFSX1 image_data_reg_34__7_ ( .D(n3087), .CK(clk), .SN(n8589), .QN(
        image_data[279]) );
  DFFSX1 image_data_reg_34__6_ ( .D(n3086), .CK(clk), .SN(n8592), .QN(
        image_data[278]) );
  DFFSX1 image_data_reg_34__5_ ( .D(n3085), .CK(clk), .SN(n8591), .QN(
        image_data[277]) );
  DFFSX1 image_data_reg_34__4_ ( .D(n3084), .CK(clk), .SN(n8590), .QN(
        image_data[276]) );
  DFFSX1 image_data_reg_34__3_ ( .D(n3083), .CK(clk), .SN(n8588), .QN(
        image_data[275]) );
  DFFSX1 image_data_reg_34__2_ ( .D(n3082), .CK(clk), .SN(n8587), .QN(
        image_data[274]) );
  DFFSX1 image_data_reg_34__1_ ( .D(n3081), .CK(clk), .SN(n8593), .QN(
        image_data[273]) );
  DFFSX1 image_data_reg_34__0_ ( .D(n3080), .CK(clk), .SN(n8576), .QN(
        image_data[272]) );
  DFFSX1 image_data_reg_33__7_ ( .D(n3079), .CK(clk), .SN(n8572), .QN(
        image_data[271]) );
  DFFSX1 image_data_reg_33__6_ ( .D(n3078), .CK(clk), .SN(n8591), .QN(
        image_data[270]) );
  DFFSX1 image_data_reg_33__5_ ( .D(n3077), .CK(clk), .SN(n8585), .QN(
        image_data[269]) );
  DFFSX1 image_data_reg_33__4_ ( .D(n3076), .CK(clk), .SN(n8576), .QN(
        image_data[268]) );
  DFFSX1 image_data_reg_33__3_ ( .D(n3075), .CK(clk), .SN(n8579), .QN(
        image_data[267]) );
  DFFSX1 image_data_reg_33__2_ ( .D(n3074), .CK(clk), .SN(n8602), .QN(
        image_data[266]) );
  DFFSX1 image_data_reg_33__1_ ( .D(n3073), .CK(clk), .SN(n8582), .QN(
        image_data[265]) );
  DFFSX1 image_data_reg_33__0_ ( .D(n3072), .CK(clk), .SN(n8598), .QN(
        image_data[264]) );
  DFFSX1 image_data_reg_32__7_ ( .D(n3071), .CK(clk), .SN(n8587), .QN(
        image_data[263]) );
  DFFSX1 image_data_reg_32__6_ ( .D(n3070), .CK(clk), .SN(n8576), .QN(
        image_data[262]) );
  DFFSX1 image_data_reg_32__5_ ( .D(n3069), .CK(clk), .SN(n8574), .QN(
        image_data[261]) );
  DFFSX1 image_data_reg_32__4_ ( .D(n3068), .CK(clk), .SN(n8571), .QN(
        image_data[260]) );
  DFFSX1 image_data_reg_32__3_ ( .D(n3067), .CK(clk), .SN(n8594), .QN(
        image_data[259]) );
  DFFSX1 image_data_reg_32__2_ ( .D(n3066), .CK(clk), .SN(n8599), .QN(
        image_data[258]) );
  DFFSX1 image_data_reg_32__1_ ( .D(n3065), .CK(clk), .SN(n8592), .QN(
        image_data[257]) );
  DFFSX1 image_data_reg_32__0_ ( .D(n3064), .CK(clk), .SN(n8597), .QN(
        image_data[256]) );
  DFFSX1 image_data_reg_31__7_ ( .D(n3063), .CK(clk), .SN(n8571), .QN(
        image_data[255]) );
  DFFSX1 image_data_reg_31__6_ ( .D(n3062), .CK(clk), .SN(n8578), .QN(
        image_data[254]) );
  DFFSX1 image_data_reg_31__5_ ( .D(n3061), .CK(clk), .SN(n8570), .QN(
        image_data[253]) );
  DFFSX1 image_data_reg_31__4_ ( .D(n3060), .CK(clk), .SN(n8581), .QN(
        image_data[252]) );
  DFFSX1 image_data_reg_31__3_ ( .D(n3059), .CK(clk), .SN(n8573), .QN(
        image_data[251]) );
  DFFSX1 image_data_reg_31__2_ ( .D(n3058), .CK(clk), .SN(n8588), .QN(
        image_data[250]) );
  DFFSX1 image_data_reg_31__1_ ( .D(n3057), .CK(clk), .SN(n8583), .QN(
        image_data[249]) );
  DFFSX1 image_data_reg_31__0_ ( .D(n3056), .CK(clk), .SN(n8571), .QN(
        image_data[248]) );
  DFFSX1 image_data_reg_30__7_ ( .D(n3055), .CK(clk), .SN(n8601), .QN(
        image_data[247]) );
  DFFSX1 image_data_reg_30__6_ ( .D(n3054), .CK(clk), .SN(n8597), .QN(
        image_data[246]) );
  DFFSX1 image_data_reg_30__5_ ( .D(n3053), .CK(clk), .SN(n8585), .QN(
        image_data[245]) );
  DFFSX1 image_data_reg_30__4_ ( .D(n3052), .CK(clk), .SN(n8584), .QN(
        image_data[244]) );
  DFFSX1 image_data_reg_30__3_ ( .D(n3051), .CK(clk), .SN(n8583), .QN(
        image_data[243]) );
  DFFSX1 image_data_reg_30__2_ ( .D(n3050), .CK(clk), .SN(n8576), .QN(
        image_data[242]) );
  DFFSX1 image_data_reg_30__1_ ( .D(n3049), .CK(clk), .SN(n8577), .QN(
        image_data[241]) );
  DFFSX1 image_data_reg_30__0_ ( .D(n3048), .CK(clk), .SN(n8578), .QN(
        image_data[240]) );
  DFFSX1 image_data_reg_29__7_ ( .D(n3047), .CK(clk), .SN(n8579), .QN(
        image_data[239]) );
  DFFSX1 image_data_reg_29__6_ ( .D(n3046), .CK(clk), .SN(n8580), .QN(
        image_data[238]) );
  DFFSX1 image_data_reg_29__5_ ( .D(n3045), .CK(clk), .SN(n8594), .QN(
        image_data[237]) );
  DFFSX1 image_data_reg_29__4_ ( .D(n3044), .CK(clk), .SN(n8595), .QN(
        image_data[236]) );
  DFFSX1 image_data_reg_29__3_ ( .D(n3043), .CK(clk), .SN(n8582), .QN(
        image_data[235]) );
  DFFSX1 image_data_reg_29__2_ ( .D(n3042), .CK(clk), .SN(n8589), .QN(
        image_data[234]) );
  DFFSX1 image_data_reg_29__1_ ( .D(n3041), .CK(clk), .SN(n8592), .QN(
        image_data[233]) );
  DFFSX1 image_data_reg_29__0_ ( .D(n3040), .CK(clk), .SN(n8591), .QN(
        image_data[232]) );
  DFFSX1 image_data_reg_28__7_ ( .D(n3039), .CK(clk), .SN(n8590), .QN(
        image_data[231]) );
  DFFSX1 image_data_reg_28__6_ ( .D(n3038), .CK(clk), .SN(n8588), .QN(
        image_data[230]) );
  DFFSX1 image_data_reg_28__5_ ( .D(n3037), .CK(clk), .SN(n8587), .QN(
        image_data[229]) );
  DFFSX1 image_data_reg_28__4_ ( .D(n3036), .CK(clk), .SN(n8593), .QN(
        image_data[228]) );
  DFFSX1 image_data_reg_28__3_ ( .D(n3035), .CK(clk), .SN(n8596), .QN(
        image_data[227]) );
  DFFSX1 image_data_reg_28__2_ ( .D(n3034), .CK(clk), .SN(n8577), .QN(
        image_data[226]) );
  DFFSX1 image_data_reg_28__1_ ( .D(n3033), .CK(clk), .SN(n8571), .QN(
        image_data[225]) );
  DFFSX1 image_data_reg_28__0_ ( .D(n3032), .CK(clk), .SN(n8576), .Q(n8560), 
        .QN(image_data[224]) );
  DFFSX1 image_data_reg_27__7_ ( .D(n3031), .CK(clk), .SN(n8585), .QN(
        image_data[223]) );
  DFFSX1 image_data_reg_27__6_ ( .D(n3030), .CK(clk), .SN(n8584), .QN(
        image_data[222]) );
  DFFSX1 image_data_reg_27__5_ ( .D(n3029), .CK(clk), .SN(n8583), .Q(n8554), 
        .QN(image_data[221]) );
  DFFSX1 image_data_reg_27__4_ ( .D(n3028), .CK(clk), .SN(n8576), .Q(n8561), 
        .QN(image_data[220]) );
  DFFSX1 image_data_reg_27__3_ ( .D(n3027), .CK(clk), .SN(n8577), .QN(
        image_data[219]) );
  DFFSX1 image_data_reg_27__2_ ( .D(n3026), .CK(clk), .SN(n8578), .QN(
        image_data[218]) );
  DFFSX1 image_data_reg_27__1_ ( .D(n3025), .CK(clk), .SN(n8579), .Q(n8562), 
        .QN(image_data[217]) );
  DFFSX1 image_data_reg_27__0_ ( .D(n3024), .CK(clk), .SN(n8580), .Q(n8555), 
        .QN(image_data[216]) );
  DFFSX1 image_data_reg_26__7_ ( .D(n3023), .CK(clk), .SN(n8594), .QN(
        image_data[215]) );
  DFFSX1 image_data_reg_26__6_ ( .D(n3022), .CK(clk), .SN(n8595), .Q(n8563), 
        .QN(image_data[214]) );
  DFFSX1 image_data_reg_26__5_ ( .D(n3021), .CK(clk), .SN(n8586), .QN(
        image_data[213]) );
  DFFSX1 image_data_reg_26__4_ ( .D(n3020), .CK(clk), .SN(n8581), .QN(
        image_data[212]) );
  DFFSX1 image_data_reg_26__3_ ( .D(n3019), .CK(clk), .SN(n8602), .QN(
        image_data[211]) );
  DFFSX1 image_data_reg_26__2_ ( .D(n3018), .CK(clk), .SN(n8575), .QN(
        image_data[210]) );
  DFFSX1 image_data_reg_26__1_ ( .D(n3017), .CK(clk), .SN(n8599), .QN(
        image_data[209]) );
  DFFSX1 image_data_reg_26__0_ ( .D(n3016), .CK(clk), .SN(n8572), .QN(
        image_data[208]) );
  DFFSX1 image_data_reg_25__7_ ( .D(n3015), .CK(clk), .SN(n8600), .QN(
        image_data[207]) );
  DFFSX1 image_data_reg_25__6_ ( .D(n3014), .CK(clk), .SN(n8573), .QN(
        image_data[206]) );
  DFFSX1 image_data_reg_25__5_ ( .D(n3013), .CK(clk), .SN(n8598), .QN(
        image_data[205]) );
  DFFSX1 image_data_reg_25__4_ ( .D(n3012), .CK(clk), .SN(n8601), .QN(
        image_data[204]) );
  DFFSX1 image_data_reg_25__3_ ( .D(n3011), .CK(clk), .SN(n8597), .QN(
        image_data[203]) );
  DFFSX1 image_data_reg_25__2_ ( .D(n3010), .CK(clk), .SN(n8585), .QN(
        image_data[202]) );
  DFFSX1 image_data_reg_25__1_ ( .D(n3009), .CK(clk), .SN(n8584), .QN(
        image_data[201]) );
  DFFSX1 image_data_reg_25__0_ ( .D(n3008), .CK(clk), .SN(n8583), .Q(n8564), 
        .QN(image_data[200]) );
  DFFSX1 image_data_reg_24__7_ ( .D(n3007), .CK(clk), .SN(n8579), .QN(
        image_data[199]) );
  DFFSX1 image_data_reg_24__6_ ( .D(n3006), .CK(clk), .SN(n8580), .QN(
        image_data[198]) );
  DFFSX1 image_data_reg_24__5_ ( .D(n3005), .CK(clk), .SN(n8594), .QN(
        image_data[197]) );
  DFFSX1 image_data_reg_24__4_ ( .D(n3004), .CK(clk), .SN(n8595), .QN(
        image_data[196]) );
  DFFSX1 image_data_reg_24__3_ ( .D(n3003), .CK(clk), .SN(n8586), .QN(
        image_data[195]) );
  DFFSX1 image_data_reg_24__2_ ( .D(n3002), .CK(clk), .SN(n8581), .QN(
        image_data[194]) );
  DFFSX1 image_data_reg_24__1_ ( .D(n3001), .CK(clk), .SN(n8582), .QN(
        image_data[193]) );
  DFFSX1 image_data_reg_24__0_ ( .D(n3000), .CK(clk), .SN(n8589), .QN(
        image_data[192]) );
  DFFSX1 image_data_reg_23__7_ ( .D(n2999), .CK(clk), .SN(n8592), .QN(
        image_data[191]) );
  DFFSX1 image_data_reg_23__6_ ( .D(n2998), .CK(clk), .SN(n8591), .QN(
        image_data[190]) );
  DFFSX1 image_data_reg_23__5_ ( .D(n2997), .CK(clk), .SN(n8590), .QN(
        image_data[189]) );
  DFFSX1 image_data_reg_23__4_ ( .D(n2996), .CK(clk), .SN(n8588), .QN(
        image_data[188]) );
  DFFSX1 image_data_reg_23__3_ ( .D(n2995), .CK(clk), .SN(n8576), .QN(
        image_data[187]) );
  DFFSX1 image_data_reg_23__2_ ( .D(n2994), .CK(clk), .SN(n8571), .QN(
        image_data[186]) );
  DFFSX1 image_data_reg_23__1_ ( .D(n2993), .CK(clk), .SN(n8583), .QN(
        image_data[185]) );
  DFFSX1 image_data_reg_23__0_ ( .D(n2992), .CK(clk), .SN(n8574), .QN(
        image_data[184]) );
  DFFSX1 image_data_reg_22__7_ ( .D(n2991), .CK(clk), .SN(n8596), .QN(
        image_data[183]) );
  DFFSX1 image_data_reg_22__6_ ( .D(n2990), .CK(clk), .SN(n8570), .QN(
        image_data[182]) );
  DFFSX1 image_data_reg_22__5_ ( .D(n2989), .CK(clk), .SN(n8602), .QN(
        image_data[181]) );
  DFFSX1 image_data_reg_22__4_ ( .D(n2988), .CK(clk), .SN(n8575), .QN(
        image_data[180]) );
  DFFSX1 image_data_reg_22__3_ ( .D(n2987), .CK(clk), .SN(n8599), .Q(n8565), 
        .QN(image_data[179]) );
  DFFSX1 image_data_reg_22__2_ ( .D(n2986), .CK(clk), .SN(n8572), .QN(
        image_data[178]) );
  DFFSX1 image_data_reg_22__1_ ( .D(n2985), .CK(clk), .SN(n8600), .QN(
        image_data[177]) );
  DFFSX1 image_data_reg_22__0_ ( .D(n2984), .CK(clk), .SN(n8573), .QN(
        image_data[176]) );
  DFFSX1 image_data_reg_21__7_ ( .D(n2983), .CK(clk), .SN(n8602), .QN(
        image_data[175]) );
  DFFSX1 image_data_reg_21__6_ ( .D(n2982), .CK(clk), .SN(n8575), .QN(
        image_data[174]) );
  DFFSX1 image_data_reg_21__5_ ( .D(n2981), .CK(clk), .SN(n8599), .QN(
        image_data[173]) );
  DFFSX1 image_data_reg_21__4_ ( .D(n2980), .CK(clk), .SN(n8572), .QN(
        image_data[172]) );
  DFFSX1 image_data_reg_21__3_ ( .D(n2979), .CK(clk), .SN(n8600), .QN(
        image_data[171]) );
  DFFSX1 image_data_reg_21__2_ ( .D(n2978), .CK(clk), .SN(n8573), .QN(
        image_data[170]) );
  DFFSX1 image_data_reg_21__1_ ( .D(n2977), .CK(clk), .SN(n8598), .QN(
        image_data[169]) );
  DFFSX1 image_data_reg_21__0_ ( .D(n2976), .CK(clk), .SN(n8601), .QN(
        image_data[168]) );
  DFFSX1 image_data_reg_20__7_ ( .D(n2975), .CK(clk), .SN(n8597), .QN(
        image_data[167]) );
  DFFSX1 image_data_reg_20__6_ ( .D(n2974), .CK(clk), .SN(n8585), .QN(
        image_data[166]) );
  DFFSX1 image_data_reg_20__5_ ( .D(n2973), .CK(clk), .SN(n8584), .QN(
        image_data[165]) );
  DFFSX1 image_data_reg_20__4_ ( .D(n2972), .CK(clk), .SN(n8583), .QN(
        image_data[164]) );
  DFFSX1 image_data_reg_20__3_ ( .D(n2971), .CK(clk), .SN(n8579), .QN(
        image_data[163]) );
  DFFSX1 image_data_reg_20__2_ ( .D(n2970), .CK(clk), .SN(n8580), .QN(
        image_data[162]) );
  DFFSX1 image_data_reg_20__1_ ( .D(n2969), .CK(clk), .SN(n8594), .QN(
        image_data[161]) );
  DFFSX1 image_data_reg_20__0_ ( .D(n2968), .CK(clk), .SN(n8595), .QN(
        image_data[160]) );
  DFFSX1 image_data_reg_19__7_ ( .D(n2967), .CK(clk), .SN(n8586), .QN(
        image_data[159]) );
  DFFSX1 image_data_reg_19__6_ ( .D(n2966), .CK(clk), .SN(n8581), .QN(
        image_data[158]) );
  DFFSX1 image_data_reg_19__5_ ( .D(n2965), .CK(clk), .SN(n8582), .QN(
        image_data[157]) );
  DFFSX1 image_data_reg_19__4_ ( .D(n2964), .CK(clk), .SN(n8589), .QN(
        image_data[156]) );
  DFFSX1 image_data_reg_19__3_ ( .D(n2963), .CK(clk), .SN(n8592), .QN(
        image_data[155]) );
  DFFSX1 image_data_reg_19__2_ ( .D(n2962), .CK(clk), .SN(n8591), .QN(
        image_data[154]) );
  DFFSX1 image_data_reg_19__1_ ( .D(n2961), .CK(clk), .SN(n8590), .QN(
        image_data[153]) );
  DFFSX1 image_data_reg_19__0_ ( .D(n2960), .CK(clk), .SN(n8588), .QN(
        image_data[152]) );
  DFFSX1 image_data_reg_18__7_ ( .D(n2959), .CK(clk), .SN(n8570), .QN(
        image_data[151]) );
  DFFSX1 image_data_reg_18__6_ ( .D(n2958), .CK(clk), .SN(n8571), .QN(
        image_data[150]) );
  DFFSX1 image_data_reg_18__5_ ( .D(n2957), .CK(clk), .SN(n8571), .QN(
        image_data[149]) );
  DFFSX1 image_data_reg_18__4_ ( .D(n2956), .CK(clk), .SN(n8577), .QN(
        image_data[148]) );
  DFFSX1 image_data_reg_18__3_ ( .D(n2955), .CK(clk), .SN(n8574), .QN(
        image_data[147]) );
  DFFSX1 image_data_reg_18__2_ ( .D(n2954), .CK(clk), .SN(n8596), .QN(
        image_data[146]) );
  DFFSX1 image_data_reg_18__1_ ( .D(n2953), .CK(clk), .SN(n8570), .QN(
        image_data[145]) );
  DFFSX1 image_data_reg_18__0_ ( .D(n2952), .CK(clk), .SN(n8602), .QN(
        image_data[144]) );
  DFFSX1 image_data_reg_17__7_ ( .D(n2951), .CK(clk), .SN(n8575), .QN(
        image_data[143]) );
  DFFSX1 image_data_reg_17__6_ ( .D(n2950), .CK(clk), .SN(n8599), .QN(
        image_data[142]) );
  DFFSX1 image_data_reg_17__5_ ( .D(n2949), .CK(clk), .SN(n8572), .QN(
        image_data[141]) );
  DFFSX1 image_data_reg_17__4_ ( .D(n2948), .CK(clk), .SN(n8600), .QN(
        image_data[140]) );
  DFFSX1 image_data_reg_17__3_ ( .D(n2947), .CK(clk), .SN(n8576), .QN(
        image_data[139]) );
  DFFSX1 image_data_reg_17__2_ ( .D(n2946), .CK(clk), .SN(n8577), .QN(
        image_data[138]) );
  DFFSX1 image_data_reg_17__1_ ( .D(n2945), .CK(clk), .SN(n8578), .QN(
        image_data[137]) );
  DFFSX1 image_data_reg_17__0_ ( .D(n2944), .CK(clk), .SN(n8579), .QN(
        image_data[136]) );
  DFFSX1 image_data_reg_16__7_ ( .D(n2943), .CK(clk), .SN(n8580), .QN(
        image_data[135]) );
  DFFSX1 image_data_reg_16__6_ ( .D(n2942), .CK(clk), .SN(n8594), .QN(
        image_data[134]) );
  DFFSX1 image_data_reg_16__5_ ( .D(n2941), .CK(clk), .SN(n8595), .QN(
        image_data[133]) );
  DFFSX1 image_data_reg_16__4_ ( .D(n2940), .CK(clk), .SN(n8586), .QN(
        image_data[132]) );
  DFFSX1 image_data_reg_16__3_ ( .D(n2939), .CK(clk), .SN(n8581), .QN(
        image_data[131]) );
  DFFSX1 image_data_reg_16__2_ ( .D(n2938), .CK(clk), .SN(n8582), .QN(
        image_data[130]) );
  DFFSX1 image_data_reg_16__1_ ( .D(n2937), .CK(clk), .SN(n8589), .QN(
        image_data[129]) );
  DFFSX1 image_data_reg_16__0_ ( .D(n2936), .CK(clk), .SN(n8592), .QN(
        image_data[128]) );
  DFFSX1 image_data_reg_15__7_ ( .D(n2935), .CK(clk), .SN(n8574), .QN(
        image_data[127]) );
  DFFSX1 image_data_reg_15__6_ ( .D(n2934), .CK(clk), .SN(n8596), .QN(
        image_data[126]) );
  DFFSX1 image_data_reg_15__5_ ( .D(n2933), .CK(clk), .SN(n8570), .QN(
        image_data[125]) );
  DFFSX1 image_data_reg_15__4_ ( .D(n2932), .CK(clk), .SN(n8602), .Q(n8547), 
        .QN(image_data[124]) );
  DFFSX1 image_data_reg_15__3_ ( .D(n2931), .CK(clk), .SN(n8575), .QN(
        image_data[123]) );
  DFFSX1 image_data_reg_15__2_ ( .D(n2930), .CK(clk), .SN(n8599), .QN(
        image_data[122]) );
  DFFSX1 image_data_reg_15__1_ ( .D(n2929), .CK(clk), .SN(n8572), .QN(
        image_data[121]) );
  DFFSX1 image_data_reg_15__0_ ( .D(n2928), .CK(clk), .SN(n8600), .QN(
        image_data[120]) );
  DFFSX1 image_data_reg_14__7_ ( .D(n2927), .CK(clk), .SN(n8573), .QN(
        image_data[119]) );
  DFFSX1 image_data_reg_14__6_ ( .D(n2926), .CK(clk), .SN(n8598), .QN(
        image_data[118]) );
  DFFSX1 image_data_reg_14__5_ ( .D(n2925), .CK(clk), .SN(n8601), .QN(
        image_data[117]) );
  DFFSX1 image_data_reg_14__4_ ( .D(n2924), .CK(clk), .SN(n8597), .QN(
        image_data[116]) );
  DFFSX1 image_data_reg_14__3_ ( .D(n2923), .CK(clk), .SN(n8590), .QN(
        image_data[115]) );
  DFFSX1 image_data_reg_14__2_ ( .D(n2922), .CK(clk), .SN(n8591), .QN(
        image_data[114]) );
  DFFSX1 image_data_reg_14__1_ ( .D(n2921), .CK(clk), .SN(n8600), .QN(
        image_data[113]) );
  DFFSX1 image_data_reg_14__0_ ( .D(n2920), .CK(clk), .SN(n8572), .QN(
        image_data[112]) );
  DFFSX1 image_data_reg_13__7_ ( .D(n2919), .CK(clk), .SN(n8571), .QN(
        image_data[111]) );
  DFFSX1 image_data_reg_13__6_ ( .D(n2918), .CK(clk), .SN(n8579), .QN(
        image_data[110]) );
  DFFSX1 image_data_reg_13__5_ ( .D(n2917), .CK(clk), .SN(n8580), .QN(
        image_data[109]) );
  DFFSX1 image_data_reg_13__4_ ( .D(n2916), .CK(clk), .SN(n8579), .QN(
        image_data[108]) );
  DFFSX1 image_data_reg_13__3_ ( .D(n2915), .CK(clk), .SN(n8575), .QN(
        image_data[107]) );
  DFFSX1 image_data_reg_13__2_ ( .D(n2914), .CK(clk), .SN(n8602), .QN(
        image_data[106]) );
  DFFSX1 image_data_reg_13__1_ ( .D(n2913), .CK(clk), .SN(n8589), .QN(
        image_data[105]) );
  DFFSX1 image_data_reg_13__0_ ( .D(n2912), .CK(clk), .SN(n8582), .QN(
        image_data[104]) );
  DFFSX1 image_data_reg_12__7_ ( .D(n2911), .CK(clk), .SN(n8599), .QN(
        image_data[103]) );
  DFFSX1 image_data_reg_12__6_ ( .D(n2910), .CK(clk), .SN(n8572), .QN(
        image_data[102]) );
  DFFSX1 image_data_reg_12__5_ ( .D(n2909), .CK(clk), .SN(n8600), .QN(
        image_data[101]) );
  DFFSX1 image_data_reg_12__4_ ( .D(n2908), .CK(clk), .SN(n8573), .QN(
        image_data[100]) );
  DFFSX1 image_data_reg_12__3_ ( .D(n2907), .CK(clk), .SN(n8598), .QN(
        image_data[99]) );
  DFFSX1 image_data_reg_12__2_ ( .D(n2906), .CK(clk), .SN(n8601), .QN(
        image_data[98]) );
  DFFSX1 image_data_reg_12__1_ ( .D(n2905), .CK(clk), .SN(n8597), .QN(
        image_data[97]) );
  DFFSX1 image_data_reg_12__0_ ( .D(n2904), .CK(clk), .SN(n8585), .QN(
        image_data[96]) );
  DFFSX1 image_data_reg_11__7_ ( .D(n2903), .CK(clk), .SN(n8584), .QN(
        image_data[95]) );
  DFFSX1 image_data_reg_11__6_ ( .D(n2902), .CK(clk), .SN(n8583), .QN(
        image_data[94]) );
  DFFSX1 image_data_reg_11__5_ ( .D(n2901), .CK(clk), .SN(n8576), .QN(
        image_data[93]) );
  DFFSX1 image_data_reg_11__4_ ( .D(n2900), .CK(clk), .SN(n8577), .QN(
        image_data[92]) );
  DFFSX1 image_data_reg_11__3_ ( .D(n2899), .CK(clk), .SN(n8599), .QN(
        image_data[91]) );
  DFFSX1 image_data_reg_11__2_ ( .D(n2898), .CK(clk), .SN(n8572), .QN(
        image_data[90]) );
  DFFSX1 image_data_reg_11__1_ ( .D(n2897), .CK(clk), .SN(n8600), .QN(
        image_data[89]) );
  DFFSX1 image_data_reg_11__0_ ( .D(n2896), .CK(clk), .SN(n8573), .QN(
        image_data[88]) );
  DFFSX1 image_data_reg_10__7_ ( .D(n2895), .CK(clk), .SN(n8598), .QN(
        image_data[87]) );
  DFFSX1 image_data_reg_10__6_ ( .D(n2894), .CK(clk), .SN(n8601), .QN(
        image_data[86]) );
  DFFSX1 image_data_reg_10__5_ ( .D(n2893), .CK(clk), .SN(n8597), .QN(
        image_data[85]) );
  DFFSX1 image_data_reg_10__4_ ( .D(n2892), .CK(clk), .SN(n8585), .QN(
        image_data[84]) );
  DFFSX1 image_data_reg_10__3_ ( .D(n2891), .CK(clk), .SN(n8584), .QN(
        image_data[83]) );
  DFFSX1 image_data_reg_10__2_ ( .D(n2890), .CK(clk), .SN(n8583), .Q(n8548), 
        .QN(image_data[82]) );
  DFFSX1 image_data_reg_10__1_ ( .D(n2889), .CK(clk), .SN(n8576), .QN(
        image_data[81]) );
  DFFSX1 image_data_reg_10__0_ ( .D(n2888), .CK(clk), .SN(n8577), .QN(
        image_data[80]) );
  DFFSX1 image_data_reg_9__7_ ( .D(n2887), .CK(clk), .SN(n8583), .QN(
        image_data[79]) );
  DFFSX1 image_data_reg_9__6_ ( .D(n2886), .CK(clk), .SN(n8574), .QN(
        image_data[78]) );
  DFFSX1 image_data_reg_9__5_ ( .D(n2885), .CK(clk), .SN(n8596), .Q(n8537), 
        .QN(image_data[77]) );
  DFFSX1 image_data_reg_9__4_ ( .D(n2884), .CK(clk), .SN(n8570), .QN(
        image_data[76]) );
  DFFSX1 image_data_reg_9__3_ ( .D(n2883), .CK(clk), .SN(n8602), .QN(
        image_data[75]) );
  DFFSX1 image_data_reg_9__2_ ( .D(n2882), .CK(clk), .SN(n8575), .Q(n8538), 
        .QN(image_data[74]) );
  DFFSX1 image_data_reg_9__1_ ( .D(n2881), .CK(clk), .SN(n8599), .QN(
        image_data[73]) );
  DFFSX1 image_data_reg_9__0_ ( .D(n2880), .CK(clk), .SN(n8572), .QN(
        image_data[72]) );
  DFFSX1 image_data_reg_8__7_ ( .D(n2879), .CK(clk), .SN(n8600), .QN(
        image_data[71]) );
  DFFSX1 image_data_reg_8__6_ ( .D(n2878), .CK(clk), .SN(n8573), .QN(
        image_data[70]) );
  DFFSX1 image_data_reg_8__5_ ( .D(n2877), .CK(clk), .SN(n8598), .QN(
        image_data[69]) );
  DFFSX1 image_data_reg_8__4_ ( .D(n2876), .CK(clk), .SN(n8601), .QN(
        image_data[68]) );
  DFFSX1 image_data_reg_8__3_ ( .D(n2875), .CK(clk), .SN(n8581), .Q(n8549), 
        .QN(image_data[67]) );
  DFFSX1 image_data_reg_8__2_ ( .D(n2874), .CK(clk), .SN(n8582), .QN(
        image_data[66]) );
  DFFSX1 image_data_reg_8__1_ ( .D(n2873), .CK(clk), .SN(n8589), .QN(
        image_data[65]) );
  DFFSX1 image_data_reg_8__0_ ( .D(n2872), .CK(clk), .SN(n8592), .QN(
        image_data[64]) );
  DFFSX1 image_data_reg_7__7_ ( .D(n2871), .CK(clk), .SN(n8591), .QN(
        image_data[63]) );
  DFFSX1 image_data_reg_7__6_ ( .D(n2870), .CK(clk), .SN(n8590), .QN(
        image_data[62]) );
  DFFSX1 image_data_reg_7__5_ ( .D(n2869), .CK(clk), .SN(n8588), .QN(
        image_data[61]) );
  DFFSX1 image_data_reg_7__4_ ( .D(n2868), .CK(clk), .SN(n8587), .QN(
        image_data[60]) );
  DFFSX1 image_data_reg_7__3_ ( .D(n2867), .CK(clk), .SN(n8593), .QN(
        image_data[59]) );
  DFFSX1 image_data_reg_7__2_ ( .D(n2866), .CK(clk), .SN(n8576), .QN(
        image_data[58]) );
  DFFSX1 image_data_reg_7__1_ ( .D(n2865), .CK(clk), .SN(n8579), .QN(
        image_data[57]) );
  DFFSX1 image_data_reg_7__0_ ( .D(n2864), .CK(clk), .SN(n8571), .QN(
        image_data[56]) );
  DFFSX1 image_data_reg_6__7_ ( .D(n2863), .CK(clk), .SN(n8588), .QN(
        image_data[55]) );
  DFFSX1 image_data_reg_6__6_ ( .D(n2862), .CK(clk), .SN(n8587), .QN(
        image_data[54]) );
  DFFSX1 image_data_reg_6__5_ ( .D(n2861), .CK(clk), .SN(n8593), .QN(
        image_data[53]) );
  DFFSX1 image_data_reg_6__4_ ( .D(n2860), .CK(clk), .SN(n8577), .QN(
        image_data[52]) );
  DFFSX1 image_data_reg_6__3_ ( .D(n2859), .CK(clk), .SN(n8583), .QN(
        image_data[51]) );
  DFFSX1 image_data_reg_6__2_ ( .D(n2858), .CK(clk), .SN(n8571), .QN(
        image_data[50]) );
  DFFSX1 image_data_reg_6__1_ ( .D(n2857), .CK(clk), .SN(n8579), .QN(
        image_data[49]) );
  DFFSX1 image_data_reg_6__0_ ( .D(n2856), .CK(clk), .SN(n8574), .QN(
        image_data[48]) );
  DFFSX1 image_data_reg_5__7_ ( .D(n2855), .CK(clk), .SN(n8596), .QN(
        image_data[47]) );
  DFFSX1 image_data_reg_5__6_ ( .D(n2854), .CK(clk), .SN(n8570), .QN(
        image_data[46]) );
  DFFSX1 image_data_reg_5__5_ ( .D(n2853), .CK(clk), .SN(n8602), .QN(
        image_data[45]) );
  DFFSX1 image_data_reg_5__4_ ( .D(n2852), .CK(clk), .SN(n8575), .QN(
        image_data[44]) );
  DFFSX1 image_data_reg_5__3_ ( .D(n2851), .CK(clk), .SN(n8594), .Q(n8550), 
        .QN(image_data[43]) );
  DFFSX1 image_data_reg_5__2_ ( .D(n2850), .CK(clk), .SN(n8595), .QN(
        image_data[42]) );
  DFFSX1 image_data_reg_5__1_ ( .D(n2849), .CK(clk), .SN(n8586), .QN(
        image_data[41]) );
  DFFSX1 image_data_reg_5__0_ ( .D(n2848), .CK(clk), .SN(n8581), .QN(
        image_data[40]) );
  DFFSX1 image_data_reg_4__7_ ( .D(n2847), .CK(clk), .SN(n8582), .QN(
        image_data[39]) );
  DFFSX1 image_data_reg_4__6_ ( .D(n2846), .CK(clk), .SN(n8589), .QN(
        image_data[38]) );
  DFFSX1 image_data_reg_4__5_ ( .D(n2845), .CK(clk), .SN(n8592), .QN(
        image_data[37]) );
  DFFSX1 image_data_reg_4__4_ ( .D(n2844), .CK(clk), .SN(n8591), .QN(
        image_data[36]) );
  DFFSX1 image_data_reg_4__3_ ( .D(n2843), .CK(clk), .SN(n8590), .QN(
        image_data[35]) );
  DFFSX1 image_data_reg_4__2_ ( .D(n2842), .CK(clk), .SN(n8588), .QN(
        image_data[34]) );
  DFFSX1 image_data_reg_4__1_ ( .D(n2841), .CK(clk), .SN(n8587), .QN(
        image_data[33]) );
  DFFSX1 image_data_reg_4__0_ ( .D(n2840), .CK(clk), .SN(n8593), .QN(
        image_data[32]) );
  DFFSX1 image_data_reg_3__7_ ( .D(n2839), .CK(clk), .SN(n8571), .QN(
        image_data[31]) );
  DFFSX1 image_data_reg_3__6_ ( .D(n2838), .CK(clk), .SN(n8574), .Q(n8551), 
        .QN(image_data[30]) );
  DFFSX1 image_data_reg_3__5_ ( .D(n2837), .CK(clk), .SN(n8596), .QN(
        image_data[29]) );
  DFFSX1 image_data_reg_3__4_ ( .D(n2836), .CK(clk), .SN(n8570), .QN(
        image_data[28]) );
  DFFSX1 image_data_reg_3__3_ ( .D(n2835), .CK(clk), .SN(n8602), .QN(
        image_data[27]) );
  DFFSX1 image_data_reg_3__2_ ( .D(n2834), .CK(clk), .SN(n8575), .QN(
        image_data[26]) );
  DFFSX1 image_data_reg_3__1_ ( .D(n2833), .CK(clk), .SN(n8599), .QN(
        image_data[25]) );
  DFFSX1 image_data_reg_3__0_ ( .D(n2832), .CK(clk), .SN(n8572), .QN(
        image_data[24]) );
  DFFSX1 image_data_reg_2__7_ ( .D(n2831), .CK(clk), .SN(n8600), .QN(
        image_data[23]) );
  DFFSX1 image_data_reg_2__6_ ( .D(n2830), .CK(clk), .SN(n8573), .QN(
        image_data[22]) );
  DFFSX1 image_data_reg_2__5_ ( .D(n2829), .CK(clk), .SN(n8598), .QN(
        image_data[21]) );
  DFFSX1 image_data_reg_2__4_ ( .D(n2828), .CK(clk), .SN(n8601), .QN(
        image_data[20]) );
  DFFSX1 image_data_reg_2__3_ ( .D(n2827), .CK(clk), .SN(n8578), .QN(
        image_data[19]) );
  DFFSX1 image_data_reg_2__2_ ( .D(n2826), .CK(clk), .SN(n8579), .QN(
        image_data[18]) );
  DFFSX1 image_data_reg_2__1_ ( .D(n2825), .CK(clk), .SN(n8580), .QN(
        image_data[17]) );
  DFFSX1 image_data_reg_2__0_ ( .D(n2824), .CK(clk), .SN(n8594), .QN(
        image_data[16]) );
  DFFSX1 image_data_reg_1__7_ ( .D(n2823), .CK(clk), .SN(n8595), .QN(
        image_data[15]) );
  DFFSX1 image_data_reg_1__6_ ( .D(n2822), .CK(clk), .SN(n8586), .QN(
        image_data[14]) );
  DFFSX1 image_data_reg_1__5_ ( .D(n2821), .CK(clk), .SN(n8581), .Q(n8552), 
        .QN(image_data[13]) );
  DFFSX1 image_data_reg_1__4_ ( .D(n2820), .CK(clk), .SN(n8582), .QN(
        image_data[12]) );
  DFFSX1 image_data_reg_1__3_ ( .D(n2819), .CK(clk), .SN(n8589), .QN(
        image_data[11]) );
  DFFSX1 image_data_reg_1__2_ ( .D(n2818), .CK(clk), .SN(n8592), .QN(
        image_data[10]) );
  DFFSX1 image_data_reg_1__1_ ( .D(n2817), .CK(clk), .SN(n8591), .QN(
        image_data[9]) );
  DFFSX1 image_data_reg_1__0_ ( .D(n2816), .CK(clk), .SN(n8590), .QN(
        image_data[8]) );
  DFFSX1 image_data_reg_0__7_ ( .D(n2815), .CK(clk), .SN(n8577), .QN(
        image_data[7]) );
  DFFSX1 image_data_reg_0__6_ ( .D(n2814), .CK(clk), .SN(n8583), .QN(
        image_data[6]) );
  DFFSX1 image_data_reg_0__5_ ( .D(n2813), .CK(clk), .SN(n8586), .QN(
        image_data[5]) );
  DFFSX1 image_data_reg_0__4_ ( .D(n2812), .CK(clk), .SN(n8573), .QN(
        image_data[4]) );
  DFFSX1 image_data_reg_0__3_ ( .D(n2811), .CK(clk), .SN(n8593), .QN(
        image_data[3]) );
  DFFSX1 image_data_reg_0__2_ ( .D(n2810), .CK(clk), .SN(n8578), .QN(
        image_data[2]) );
  DFFSX1 image_data_reg_0__1_ ( .D(n2809), .CK(clk), .SN(n8581), .QN(
        image_data[1]) );
  DFFSX1 image_data_reg_0__0_ ( .D(n2808), .CK(clk), .SN(n8598), .QN(
        image_data[0]) );
  CMPR42X1 DP_OP_2677J1_122_9848_U16 ( .A(n8569), .B(N2760), .C(N2784), .D(
        N2776), .ICI(DP_OP_2677J1_122_9848_n30), .S(DP_OP_2677J1_122_9848_n27), 
        .ICO(DP_OP_2677J1_122_9848_n25), .CO(DP_OP_2677J1_122_9848_n26) );
  CMPR42X1 DP_OP_2677J1_122_9848_U15 ( .A(n8568), .B(N2759), .C(N2783), .D(
        N2775), .ICI(DP_OP_2677J1_122_9848_n25), .S(DP_OP_2677J1_122_9848_n24), 
        .ICO(DP_OP_2677J1_122_9848_n22), .CO(DP_OP_2677J1_122_9848_n23) );
  CMPR42X1 DP_OP_2677J1_122_9848_U14 ( .A(N2766), .B(N2758), .C(N2782), .D(
        N2774), .ICI(DP_OP_2677J1_122_9848_n22), .S(DP_OP_2677J1_122_9848_n21), 
        .ICO(DP_OP_2677J1_122_9848_n19), .CO(DP_OP_2677J1_122_9848_n20) );
  CMPR42X1 DP_OP_2677J1_122_9848_U13 ( .A(N2765), .B(N2757), .C(N2781), .D(
        N2773), .ICI(DP_OP_2677J1_122_9848_n19), .S(DP_OP_2677J1_122_9848_n18), 
        .ICO(DP_OP_2677J1_122_9848_n16), .CO(DP_OP_2677J1_122_9848_n17) );
  CMPR42X1 DP_OP_2677J1_122_9848_U12 ( .A(n8567), .B(N2756), .C(N2780), .D(
        N2772), .ICI(DP_OP_2677J1_122_9848_n16), .S(DP_OP_2677J1_122_9848_n15), 
        .ICO(DP_OP_2677J1_122_9848_n13), .CO(DP_OP_2677J1_122_9848_n14) );
  CMPR42X1 DP_OP_2677J1_122_9848_U11 ( .A(n3442), .B(N2755), .C(N2779), .D(
        N2771), .ICI(DP_OP_2677J1_122_9848_n13), .S(DP_OP_2677J1_122_9848_n12), 
        .ICO(DP_OP_2677J1_122_9848_n10), .CO(DP_OP_2677J1_122_9848_n11) );
  DFFSX1 IROM_rd_reg ( .D(n3340), .CK(clk), .SN(n8580), .Q(IROM_rd), .QN(n8566) );
  DFFSX1 busy_reg ( .D(n3343), .CK(clk), .SN(n8596), .Q(busy), .QN(n8534) );
  DFFSX1 cs_reg_1_ ( .D(n3327), .CK(clk), .SN(n8581), .Q(n8533), .QN(cs[1]) );
  DFFSX1 IRAM_valid_reg ( .D(n3320), .CK(clk), .SN(n8591), .QN(IRAM_valid) );
  DFFSX1 out_done_reg ( .D(n3339), .CK(clk), .SN(n8582), .QN(done) );
  DFFSX1 cs_reg_0_ ( .D(n3328), .CK(clk), .SN(n8589), .QN(cs[0]) );
  DFFSX4 y_pos_reg_2_ ( .D(n3330), .CK(clk), .SN(n8571), .Q(n8521), .QN(
        IROM_A[5]) );
  DFFSX2 x_pos_reg_2_ ( .D(n3332), .CK(clk), .SN(n8583), .Q(n8519), .QN(
        IROM_A[2]) );
  DFFSX2 y_cal_reg_2_ ( .D(n3342), .CK(clk), .SN(n8576), .Q(op4[5]), .QN(n8525) );
  DFFSX2 y_cal_reg_0_ ( .D(n3326), .CK(clk), .SN(n8578), .Q(n8524), .QN(op4[3]) );
  DFFSX2 x_pos_reg_0_ ( .D(n3333), .CK(clk), .SN(n8578), .Q(n8526), .QN(
        IROM_A[0]) );
  DFFSX2 x_pos_reg_1_ ( .D(n3338), .CK(clk), .SN(n8577), .Q(n8520), .QN(
        IROM_A[1]) );
  DFFSX2 y_pos_reg_0_ ( .D(n3321), .CK(clk), .SN(n8595), .Q(n8522), .QN(
        IROM_A[3]) );
  DFFSX2 y_pos_reg_1_ ( .D(n3331), .CK(clk), .SN(n8579), .Q(n8527), .QN(
        IROM_A[4]) );
  DFFSX2 x_cal_reg_2_ ( .D(n3341), .CK(clk), .SN(n8574), .Q(op2[2]), .QN(n8528) );
  DFFSX1 x_cal_reg_0_ ( .D(n3324), .CK(clk), .SN(n8595), .Q(n8529), .QN(op2[0]) );
  AOI211X1 U3373 ( .A0(n8333), .A1(n3352), .B0(n6887), .C0(n6886), .Y(n3278)
         );
  AOI211X1 U3374 ( .A0(n8503), .A1(n8333), .B0(n6866), .C0(n6865), .Y(n3276)
         );
  AOI211X1 U3375 ( .A0(n3351), .A1(n8333), .B0(n6933), .C0(n6932), .Y(n3273)
         );
  AOI211X1 U3376 ( .A0(n3369), .A1(n8333), .B0(n8332), .C0(n8331), .Y(n3275)
         );
  AOI211X1 U3377 ( .A0(n3362), .A1(n8333), .B0(n6914), .C0(n6913), .Y(n3279)
         );
  INVX4 U3378 ( .A(n3385), .Y(n3356) );
  INVX4 U3379 ( .A(n3386), .Y(n3349) );
  INVX1 U3380 ( .A(n7303), .Y(n3464) );
  CLKINVX3 U3381 ( .A(n6951), .Y(n3392) );
  INVX1 U3382 ( .A(n6893), .Y(n6787) );
  INVX1 U3383 ( .A(n8430), .Y(n8454) );
  NOR4X1 U3384 ( .A(n3905), .B(n3904), .C(n3903), .D(n3902), .Y(n3927) );
  NOR4XL U3385 ( .A(n3925), .B(n3924), .C(n3923), .D(n3922), .Y(n3926) );
  BUFX1 U3386 ( .A(n6919), .Y(n3437) );
  CLKINVX3 U3387 ( .A(n6973), .Y(n3393) );
  INVX4 U3388 ( .A(n3396), .Y(n3350) );
  INVX4 U3389 ( .A(n3419), .Y(n3360) );
  CLKINVX8 U3390 ( .A(n3418), .Y(n6855) );
  CLKINVX3 U3391 ( .A(n3440), .Y(n3365) );
  INVX4 U3392 ( .A(n3439), .Y(n3344) );
  INVX4 U3393 ( .A(n3440), .Y(n3345) );
  INVX4 U3394 ( .A(n3437), .Y(n3346) );
  INVX8 U3395 ( .A(n6403), .Y(n3347) );
  CLKINVX8 U3396 ( .A(n6827), .Y(n3348) );
  CLKBUFX3 U3397 ( .A(n5025), .Y(n3462) );
  CLKBUFX3 U3398 ( .A(n5209), .Y(n3460) );
  CLKBUFX3 U3399 ( .A(n5037), .Y(n3458) );
  BUFX3 U3400 ( .A(n5197), .Y(n3463) );
  CLKBUFX3 U3401 ( .A(n5051), .Y(n3457) );
  CLKBUFX3 U3402 ( .A(n5223), .Y(n3459) );
  NAND2X1 U3403 ( .A(n5004), .B(n5171), .Y(n5003) );
  NAND2X1 U3404 ( .A(n5173), .B(n5171), .Y(n5172) );
  CLKINVX3 U3405 ( .A(n3394), .Y(n3368) );
  INVX4 U3406 ( .A(n8199), .Y(n3369) );
  CLKINVX4 U3407 ( .A(n6787), .Y(n3394) );
  CLKINVX4 U3408 ( .A(n3370), .Y(n3388) );
  AOI2BB2XL U3409 ( .B0(n8114), .B1(n3382), .A0N(n3397), .A1N(n3419), .Y(n6988) );
  BUFX2 U3410 ( .A(n7035), .Y(n6651) );
  CLKINVX4 U3411 ( .A(n3390), .Y(n3373) );
  BUFX2 U3412 ( .A(n8341), .Y(n6291) );
  BUFX2 U3413 ( .A(n7690), .Y(n7581) );
  CLKINVX4 U3414 ( .A(n6852), .Y(n3370) );
  CLKINVX3 U3415 ( .A(n7761), .Y(n3372) );
  BUFX2 U3416 ( .A(n7487), .Y(n7326) );
  BUFX2 U3417 ( .A(n7902), .Y(n6880) );
  INVX8 U3418 ( .A(n7980), .Y(n3351) );
  INVX8 U3419 ( .A(n8509), .Y(n3352) );
  INVXL U3420 ( .A(n8340), .Y(n8372) );
  CLKINVX8 U3421 ( .A(n3392), .Y(n3353) );
  INVX2 U3422 ( .A(n7191), .Y(n3374) );
  CLKINVX8 U3423 ( .A(n3393), .Y(n3354) );
  NOR2X1 U3424 ( .A(n3454), .B(n6998), .Y(n8031) );
  BUFX2 U3425 ( .A(n7261), .Y(n6979) );
  INVX4 U3426 ( .A(n3390), .Y(n3355) );
  BUFX2 U3427 ( .A(n7930), .Y(n7078) );
  CLKINVX8 U3428 ( .A(n3391), .Y(n3357) );
  BUFX3 U3429 ( .A(n6879), .Y(n7795) );
  OR2X2 U3430 ( .A(n6176), .B(n6583), .Y(n6407) );
  INVX4 U3431 ( .A(n7773), .Y(n3358) );
  CLKINVX3 U3432 ( .A(n3375), .Y(n3359) );
  INVX8 U3433 ( .A(n7307), .Y(n3361) );
  INVX8 U3434 ( .A(n7578), .Y(n3362) );
  INVX1 U3435 ( .A(N2773), .Y(n4971) );
  AOI22X2 U3436 ( .A0(n5168), .A1(n3927), .B0(n3926), .B1(n4868), .Y(N2776) );
  NOR4X1 U3437 ( .A(n3599), .B(n3598), .C(n3597), .D(n3596), .Y(n3600) );
  NOR4X1 U3438 ( .A(n4169), .B(n4168), .C(n4167), .D(n4166), .Y(n4191) );
  NOR4XL U3439 ( .A(n4490), .B(n4489), .C(n4488), .D(n4487), .Y(n4491) );
  NOR4X1 U3440 ( .A(n4189), .B(n4188), .C(n4187), .D(n4186), .Y(n4190) );
  NOR4XL U3441 ( .A(n4470), .B(n4469), .C(n4468), .D(n4467), .Y(n4492) );
  NOR4X1 U3442 ( .A(n3579), .B(n3578), .C(n3577), .D(n3576), .Y(n3601) );
  CLKBUFX2 U3443 ( .A(n8280), .Y(n3452) );
  NOR2X4 U3444 ( .A(n8524), .B(n8500), .Y(n5908) );
  OR2XL U3445 ( .A(n6401), .B(n6758), .Y(n6341) );
  OR2X1 U3446 ( .A(n7029), .B(n6767), .Y(n4589) );
  CLKINVX8 U3447 ( .A(n3398), .Y(n3363) );
  OR2XL U3448 ( .A(n7029), .B(n6710), .Y(n5924) );
  BUFX2 U3449 ( .A(n8491), .Y(n3451) );
  OR2XL U3450 ( .A(n6747), .B(n7029), .Y(n8500) );
  BUFX3 U3451 ( .A(n4768), .Y(n3896) );
  CLKINVX8 U3452 ( .A(n5010), .Y(n3364) );
  BUFX3 U3453 ( .A(n3791), .Y(n3928) );
  BUFX3 U3454 ( .A(n4670), .Y(n3897) );
  OR2XL U3455 ( .A(n8483), .B(n6766), .Y(n5707) );
  BUFX3 U3456 ( .A(n3798), .Y(n3887) );
  BUFX3 U3457 ( .A(n4428), .Y(n3936) );
  BUFX3 U3458 ( .A(n4753), .Y(n3865) );
  BUFX3 U3459 ( .A(n4433), .Y(n3941) );
  BUFX3 U3460 ( .A(n4713), .Y(n3866) );
  BUFX3 U3461 ( .A(n3804), .Y(n3867) );
  BUFX3 U3462 ( .A(n4754), .Y(n3942) );
  BUFX3 U3463 ( .A(n3797), .Y(n3886) );
  BUFX3 U3464 ( .A(n4434), .Y(n3943) );
  BUFX3 U3465 ( .A(n4720), .Y(n3874) );
  BUFX3 U3466 ( .A(n4439), .Y(n3948) );
  BUFX3 U3467 ( .A(n3810), .Y(n3876) );
  OR2XL U3468 ( .A(n6748), .B(n6726), .Y(n8349) );
  BUFX3 U3469 ( .A(n4722), .Y(n3877) );
  BUFX3 U3470 ( .A(n4440), .Y(n3949) );
  BUFX3 U3471 ( .A(n4708), .Y(n3884) );
  BUFX3 U3472 ( .A(n4422), .Y(n3929) );
  BUFX3 U3473 ( .A(n3792), .Y(n3894) );
  BUFX3 U3474 ( .A(n4427), .Y(n3934) );
  BUFX3 U3475 ( .A(n3805), .Y(n3869) );
  OR2XL U3476 ( .A(n7034), .B(n6710), .Y(n6146) );
  OR2XL U3477 ( .A(n3438), .B(n6766), .Y(n6290) );
  BUFX3 U3478 ( .A(n3811), .Y(n3879) );
  BUFX3 U3479 ( .A(n3799), .Y(n3888) );
  NOR2X4 U3480 ( .A(n8519), .B(n8489), .Y(IRAM_A[2]) );
  INVX1 U3481 ( .A(n4595), .Y(n5255) );
  NAND2XL U3482 ( .A(n8518), .B(op4[5]), .Y(n6747) );
  NOR2X1 U3483 ( .A(op2[2]), .B(op4[3]), .Y(n3470) );
  AOI221XL U3484 ( .A0(image_data[72]), .A1(n3454), .B0(n7001), .B1(n8018), 
        .C0(n7000), .Y(n2880) );
  AOI211XL U3485 ( .A0(n3352), .A1(n8348), .B0(n7726), .C0(n7725), .Y(n3270)
         );
  BUFX3 U3486 ( .A(n6586), .Y(n6959) );
  AOI32XL U3487 ( .A0(n3348), .A1(n8018), .A2(n6947), .B0(n8028), .B1(n8538), 
        .Y(n6948) );
  CLKINVX3 U3488 ( .A(n6585), .Y(n6586) );
  CLKINVX4 U3489 ( .A(n3437), .Y(n3366) );
  CLKINVX4 U3490 ( .A(n3439), .Y(n3367) );
  BUFX3 U3491 ( .A(n6854), .Y(n3418) );
  OAI21XL U3492 ( .A0(n6020), .A1(n6583), .B0(n6019), .Y(n6837) );
  AOI222X1 U3493 ( .A0(n6581), .A1(n5797), .B0(n6579), .B1(n5796), .C0(n6577), 
        .C1(n5795), .Y(n5799) );
  AOI222X1 U3494 ( .A0(n6581), .A1(n6580), .B0(n6579), .B1(n6578), .C0(n6577), 
        .C1(n6576), .Y(n6584) );
  AOI222X1 U3495 ( .A0(n6581), .A1(n6120), .B0(n6579), .B1(n6119), .C0(n6577), 
        .C1(n6118), .Y(n6122) );
  AOI222X1 U3496 ( .A0(n6581), .A1(n5695), .B0(n6579), .B1(n5694), .C0(n6577), 
        .C1(n5693), .Y(n5697) );
  AOI222X1 U3497 ( .A0(n6581), .A1(n5900), .B0(n6579), .B1(n5899), .C0(n6577), 
        .C1(n5898), .Y(n5902) );
  BUFX2 U3498 ( .A(n5203), .Y(n3448) );
  BUFX2 U3499 ( .A(n5031), .Y(n3447) );
  INVX1 U3500 ( .A(n5043), .Y(n5030) );
  INVX1 U3501 ( .A(n5215), .Y(n5202) );
  NAND2BX1 U3502 ( .AN(n4997), .B(n4998), .Y(n5008) );
  NAND2X1 U3503 ( .A(n5164), .B(n5163), .Y(n5179) );
  NOR2X1 U3504 ( .A(n5185), .B(n5166), .Y(n5164) );
  BUFX2 U3505 ( .A(n6943), .Y(n6332) );
  CLKINVX3 U3506 ( .A(n8372), .Y(n3387) );
  INVX2 U3507 ( .A(n7773), .Y(n7923) );
  CLKINVX8 U3508 ( .A(n8035), .Y(n3371) );
  NAND2X1 U3509 ( .A(n4978), .B(n3442), .Y(n5160) );
  AOI22X1 U3510 ( .A0(N2776), .A1(n6421), .B0(n8569), .B1(n6420), .Y(n7754) );
  OR2X2 U3511 ( .A(n5269), .B(n6583), .Y(n7773) );
  CLKINVX8 U3512 ( .A(n7068), .Y(n3375) );
  CLKINVX2 U3513 ( .A(n8084), .Y(n8185) );
  AOI22X2 U3514 ( .A0(op4[5]), .A1(n4637), .B0(n4636), .B1(n8525), .Y(n6126)
         );
  AOI22X2 U3515 ( .A0(op4[5]), .A1(n4191), .B0(n4190), .B1(n8525), .Y(N2766)
         );
  OAI221X4 U3516 ( .A0(in_valid), .A1(IRAM_D[2]), .B0(n8523), .B1(IROM_Q[2]), 
        .C0(n8480), .Y(n5266) );
  OAI221X4 U3517 ( .A0(in_valid), .A1(IRAM_D[3]), .B0(n8523), .B1(IROM_Q[3]), 
        .C0(n8480), .Y(n6265) );
  NOR4X1 U3518 ( .A(n4399), .B(n4398), .C(n4397), .D(n4396), .Y(n4400) );
  NOR4X1 U3519 ( .A(n4379), .B(n4378), .C(n4377), .D(n4376), .Y(n4401) );
  INVX4 U3520 ( .A(n5168), .Y(n4868) );
  AOI22XL U3521 ( .A0(n6779), .A1(n6904), .B0(n3398), .B1(n6398), .Y(n6963) );
  CLKINVX2 U3522 ( .A(n8385), .Y(n7995) );
  CLKINVX4 U3523 ( .A(n6352), .Y(n3376) );
  CLKINVX2 U3524 ( .A(n8200), .Y(n8393) );
  BUFX3 U3525 ( .A(n4681), .Y(n3895) );
  CLKINVX4 U3526 ( .A(n5924), .Y(n3377) );
  CLKINVX2 U3527 ( .A(n8125), .Y(n8490) );
  CLKINVX4 U3528 ( .A(n6341), .Y(n3378) );
  AND2XL U3529 ( .A(n6639), .B(n6992), .Y(n6641) );
  CLKINVX4 U3530 ( .A(n4589), .Y(n3379) );
  CLKINVX4 U3531 ( .A(n6165), .Y(n3380) );
  CLKINVX4 U3532 ( .A(n5907), .Y(n3381) );
  BUFX3 U3533 ( .A(n4714), .Y(n3868) );
  BUFX3 U3534 ( .A(n4707), .Y(n3885) );
  CLKINVX4 U3535 ( .A(n5707), .Y(n3382) );
  BUFX3 U3536 ( .A(n4702), .Y(n3893) );
  BUFX3 U3537 ( .A(n4721), .Y(n3878) );
  BUFX3 U3538 ( .A(n4719), .Y(n3875) );
  BUFX3 U3539 ( .A(n4763), .Y(n3935) );
  OR2XL U3540 ( .A(n6742), .B(n6792), .Y(n6398) );
  NOR2X4 U3541 ( .A(n5002), .B(n3482), .Y(n4681) );
  CLKINVX4 U3542 ( .A(n6146), .Y(n3383) );
  NOR2X2 U3543 ( .A(n6384), .B(n5255), .Y(n6581) );
  CLKINVX4 U3544 ( .A(n6290), .Y(n3384) );
  BUFX2 U3545 ( .A(n4555), .Y(n3456) );
  NOR2XL U3546 ( .A(cmd_reg[3]), .B(n8532), .Y(n4595) );
  NOR2XL U3547 ( .A(cmd_reg[1]), .B(n8531), .Y(n6303) );
  INVX8 U3548 ( .A(n8524), .Y(n6401) );
  NAND2X1 U3549 ( .A(n8531), .B(cmd_reg[1]), .Y(n6304) );
  AOI211XL U3550 ( .A0(n8503), .A1(n8339), .B0(n7516), .C0(n7515), .Y(n3244)
         );
  AOI211XL U3551 ( .A0(n8503), .A1(n8286), .B0(n7443), .C0(n7442), .Y(n3228)
         );
  AOI211XL U3552 ( .A0(n3373), .A1(n8348), .B0(n7520), .C0(n7519), .Y(n3264)
         );
  AOI211XL U3553 ( .A0(n8079), .A1(image_data[448]), .B0(n8078), .C0(n8077), 
        .Y(n3256) );
  AOI211XL U3554 ( .A0(n3373), .A1(n8333), .B0(n6815), .C0(n6814), .Y(n3272)
         );
  AOI211XL U3555 ( .A0(n3355), .A1(n8436), .B0(n8113), .C0(n8112), .Y(n2856)
         );
  AOI211XL U3556 ( .A0(n3454), .A1(image_data[78]), .B0(n7585), .C0(n7584), 
        .Y(n2886) );
  AOI211XL U3557 ( .A0(n8503), .A1(n7486), .B0(n6394), .C0(n6393), .Y(n3108)
         );
  AOI211XL U3558 ( .A0(n3373), .A1(n8286), .B0(n7457), .C0(n7456), .Y(n3224)
         );
  AOI211XL U3559 ( .A0(n3373), .A1(n8339), .B0(n7512), .C0(n7511), .Y(n3240)
         );
  AOI211XL U3560 ( .A0(n8259), .A1(n7078), .B0(n3464), .C0(n6336), .Y(n6339)
         );
  AOI211XL U3561 ( .A0(n3380), .A1(n6979), .B0(n3464), .C0(n6342), .Y(n6344)
         );
  AOI211XL U3562 ( .A0(n3369), .A1(n8436), .B0(n8435), .C0(n8434), .Y(n2859)
         );
  AOI211XL U3563 ( .A0(n7795), .A1(n7486), .B0(n6397), .C0(n6396), .Y(n3106)
         );
  AOI32XL U3564 ( .A0(n7303), .A1(n8018), .A2(n7055), .B0(n8028), .B1(n8537), 
        .Y(n7056) );
  BUFX3 U3565 ( .A(n6810), .Y(n3439) );
  BUFX3 U3566 ( .A(n6797), .Y(n3440) );
  CLKINVX4 U3567 ( .A(n6837), .Y(n7303) );
  AOI222X4 U3568 ( .A0(n6581), .A1(n5265), .B0(n6579), .B1(n5264), .C0(n6577), 
        .C1(n5263), .Y(n5267) );
  AOI222X4 U3569 ( .A0(n6581), .A1(n6264), .B0(n6579), .B1(n6263), .C0(n6577), 
        .C1(n6262), .Y(n6266) );
  INVX1 U3570 ( .A(n6498), .Y(n6495) );
  AOI22XL U3571 ( .A0(op2[0]), .A1(n5173), .B0(n5175), .B1(n8529), .Y(n5215)
         );
  INVX1 U3572 ( .A(n6574), .Y(n6571) );
  AOI22XL U3573 ( .A0(op2[0]), .A1(n5004), .B0(n5005), .B1(n8529), .Y(n5043)
         );
  INVX2 U3574 ( .A(n5005), .Y(n5004) );
  INVX2 U3575 ( .A(n5175), .Y(n5173) );
  INVX1 U3576 ( .A(n5008), .Y(n5012) );
  NOR2XL U3577 ( .A(n5015), .B(n4999), .Y(n4998) );
  NAND4BXL U3578 ( .AN(n5125), .B(n5124), .C(n5123), .D(n5122), .Y(n5177) );
  AND4XL U3579 ( .A(n5149), .B(n5148), .C(n5147), .D(n5146), .Y(n5166) );
  OAI32XL U3580 ( .A0(n8501), .A1(n6786), .A2(n8199), .B0(n8447), .B1(n7907), 
        .Y(n6373) );
  AOI2BB1XL U3581 ( .A0N(n5091), .A1N(n5090), .B0(n5089), .Y(n5094) );
  CLKBUFX3 U3582 ( .A(n7507), .Y(n3419) );
  INVX4 U3583 ( .A(n7517), .Y(n3385) );
  CLKINVX8 U3584 ( .A(n8111), .Y(n8114) );
  INVX2 U3585 ( .A(n6407), .Y(n8423) );
  AND2XL U3586 ( .A(n5910), .B(n8160), .Y(n8163) );
  CLKINVX4 U3587 ( .A(n8376), .Y(n3386) );
  AND2XL U3588 ( .A(n5923), .B(n8178), .Y(n8181) );
  CLKINVX4 U3589 ( .A(n6407), .Y(n3389) );
  INVX2 U3590 ( .A(n6346), .Y(n3390) );
  AND3XL U3591 ( .A(n8446), .B(n6795), .C(n8250), .Y(n8253) );
  AND3XL U3592 ( .A(n8406), .B(n8400), .C(n7010), .Y(n8403) );
  AND3XL U3593 ( .A(n8432), .B(n6824), .C(n8245), .Y(n8248) );
  INVX4 U3594 ( .A(n7938), .Y(n3391) );
  INVX4 U3595 ( .A(n7754), .Y(n3395) );
  CLKINVX4 U3596 ( .A(n7723), .Y(n3396) );
  INVXL U3597 ( .A(N2760), .Y(n4986) );
  INVXL U3598 ( .A(N2782), .Y(n5704) );
  INVXL U3599 ( .A(N2776), .Y(n4966) );
  AND2XL U3600 ( .A(n6160), .B(n8172), .Y(n8175) );
  INVXL U3601 ( .A(N2775), .Y(n4967) );
  INVXL U3602 ( .A(N2780), .Y(n5807) );
  INVXL U3603 ( .A(n8459), .Y(n4985) );
  INVX2 U3604 ( .A(n7009), .Y(n8400) );
  INVXL U3605 ( .A(N2755), .Y(n4993) );
  INVXL U3606 ( .A(N2774), .Y(n4964) );
  AND2XL U3607 ( .A(n6167), .B(n8166), .Y(n8169) );
  INVXL U3608 ( .A(N2765), .Y(n4989) );
  INVX2 U3609 ( .A(n6823), .Y(n8245) );
  INVX2 U3610 ( .A(n6794), .Y(n8250) );
  AND2XL U3611 ( .A(n6592), .B(n8137), .Y(n8140) );
  INVXL U3612 ( .A(n8458), .Y(n5603) );
  AOI22X2 U3613 ( .A0(n5168), .A1(n4870), .B0(n4869), .B1(n4868), .Y(n4871) );
  INVX2 U3614 ( .A(n3441), .Y(n3442) );
  AND2XL U3615 ( .A(n7983), .B(n8143), .Y(n8146) );
  AOI22X2 U3616 ( .A0(n3450), .A1(n4492), .B0(n4491), .B1(n4959), .Y(N2758) );
  AND2XL U3617 ( .A(n5709), .B(n8394), .Y(n8397) );
  BUFX2 U3618 ( .A(n3728), .Y(n8567) );
  NOR4XL U3619 ( .A(n4042), .B(n4041), .C(n4040), .D(n4039), .Y(n4064) );
  AND2XL U3620 ( .A(n7972), .B(n8154), .Y(n8157) );
  NOR4XL U3621 ( .A(n3537), .B(n3536), .C(n3535), .D(n3534), .Y(n3559) );
  INVX1 U3622 ( .A(N2763), .Y(n3441) );
  AND3XL U3623 ( .A(n8310), .B(n6348), .C(n8240), .Y(n8243) );
  INVXL U3624 ( .A(N2766), .Y(n4990) );
  AND3XL U3625 ( .A(n6668), .B(n7684), .C(n8203), .Y(n8206) );
  NOR4XL U3626 ( .A(n4062), .B(n4061), .C(n4060), .D(n4059), .Y(n4063) );
  AND3XL U3627 ( .A(n6616), .B(n8209), .C(n8195), .Y(n8198) );
  AND3XL U3628 ( .A(n8159), .B(n6658), .C(n8230), .Y(n8233) );
  AND3XL U3629 ( .A(n6634), .B(n8289), .C(n8190), .Y(n8193) );
  NOR4XL U3630 ( .A(n3557), .B(n3556), .C(n3555), .D(n3554), .Y(n3558) );
  AOI22X2 U3631 ( .A0(n5168), .A1(n4401), .B0(n4400), .B1(n4868), .Y(N2771) );
  INVX2 U3632 ( .A(n6657), .Y(n8230) );
  INVX2 U3633 ( .A(n6649), .Y(n8218) );
  INVX2 U3634 ( .A(n6615), .Y(n8195) );
  INVX2 U3635 ( .A(n6633), .Y(n8190) );
  AOI21XL U3636 ( .A0(n7032), .A1(n6779), .B0(n6356), .Y(n6978) );
  INVX2 U3637 ( .A(n6667), .Y(n8203) );
  INVX2 U3638 ( .A(n7907), .Y(n8501) );
  NOR4XL U3639 ( .A(n3495), .B(n3494), .C(n3493), .D(n3492), .Y(n3517) );
  AND3XL U3640 ( .A(n6627), .B(n8304), .C(n8210), .Y(n8213) );
  NOR4XL U3641 ( .A(n3515), .B(n3514), .C(n3513), .D(n3512), .Y(n3516) );
  NOR2XL U3642 ( .A(n7043), .B(n7042), .Y(n7046) );
  INVX2 U3643 ( .A(n8165), .Y(n8238) );
  INVX2 U3644 ( .A(n6626), .Y(n8210) );
  BUFX3 U3645 ( .A(n5167), .Y(n3450) );
  INVX2 U3646 ( .A(n8159), .Y(n8228) );
  OR2XL U3647 ( .A(n6802), .B(n6777), .Y(n6352) );
  INVXL U3648 ( .A(n8446), .Y(n8032) );
  INVX2 U3649 ( .A(n8370), .Y(n8182) );
  INVX2 U3650 ( .A(n8215), .Y(n8310) );
  CLKINVX4 U3651 ( .A(n6641), .Y(n3397) );
  OR2XL U3652 ( .A(n8524), .B(n6634), .Y(n5907) );
  INVX2 U3653 ( .A(n8406), .Y(n8398) );
  OR2XL U3654 ( .A(n8524), .B(n6758), .Y(n6165) );
  INVX1 U3655 ( .A(n8467), .Y(n5009) );
  INVX2 U3656 ( .A(n8136), .Y(n7888) );
  CLKINVX3 U3657 ( .A(n6337), .Y(n3398) );
  NAND2X2 U3658 ( .A(n3449), .B(n5929), .Y(n3399) );
  INVX2 U3659 ( .A(n3405), .Y(n8342) );
  NOR2X4 U3660 ( .A(n6374), .B(n6401), .Y(n6143) );
  AOI31XL U3661 ( .A0(cs[0]), .A1(n8533), .A2(n8461), .B0(n8488), .Y(n8462) );
  AOI31XL U3662 ( .A0(cs[0]), .A1(cmd_valid), .A2(n8461), .B0(n8460), .Y(n6323) );
  NOR2X2 U3663 ( .A(n5255), .B(n6310), .Y(n6577) );
  NAND2XL U3664 ( .A(op4[3]), .B(n6991), .Y(n6726) );
  NOR2X2 U3665 ( .A(n5255), .B(n6304), .Y(n6579) );
  AND2XL U3666 ( .A(n8480), .B(n8481), .Y(n7043) );
  NOR3BXL U3667 ( .AN(n7040), .B(n8527), .C(n7039), .Y(n8481) );
  INVX2 U3668 ( .A(n3400), .Y(n3438) );
  CLKINVX4 U3669 ( .A(n4590), .Y(n6583) );
  NAND2X2 U3670 ( .A(op2[1]), .B(n8529), .Y(n3471) );
  NOR3X2 U3671 ( .A(IROM_A[0]), .B(n8520), .C(n8519), .Y(n3410) );
  OR4XL U3672 ( .A(cmd[0]), .B(cmd[1]), .C(cmd[2]), .D(cmd[3]), .Y(n8461) );
  OAI22XL U3673 ( .A0(n4871), .A1(n5604), .B0(N2776), .B1(n4872), .Y(n5109) );
  INVXL U3674 ( .A(n6127), .Y(n5098) );
  AOI21XL U3675 ( .A0(N2782), .A1(n4964), .B0(n4874), .Y(n5112) );
  NAND2XL U3676 ( .A(N2781), .B(n4971), .Y(n4873) );
  OAI22XL U3677 ( .A0(N2783), .A1(n4967), .B0(N2784), .B1(n4966), .Y(n5113) );
  OAI22XL U3678 ( .A0(N2784), .A1(n4986), .B0(n5698), .B1(n5603), .Y(n5127) );
  AOI22XL U3679 ( .A0(N2784), .A1(n4986), .B0(N2783), .B1(n6173), .Y(n5126) );
  AOI22XL U3680 ( .A0(N2757), .A1(n4971), .B0(N2756), .B1(n5115), .Y(n5092) );
  OAI22XL U3681 ( .A0(N2757), .A1(n4971), .B0(N2758), .B1(n4964), .Y(n5093) );
  AOI22XL U3682 ( .A0(N2774), .A1(n4990), .B0(N2775), .B1(n4984), .Y(n5105) );
  OAI22XL U3683 ( .A0(N2774), .A1(n4990), .B0(N2773), .B1(n4989), .Y(n5103) );
  NAND2XL U3684 ( .A(n8459), .B(n5604), .Y(n5150) );
  NAND3BXL U3685 ( .AN(n6126), .B(n6123), .C(n5150), .Y(n5153) );
  AOI22XL U3686 ( .A0(N2758), .A1(n4990), .B0(N2759), .B1(n4984), .Y(n5142) );
  OAI22XL U3687 ( .A0(N2758), .A1(n4990), .B0(N2757), .B1(n4989), .Y(n5140) );
  AOI21XL U3688 ( .A0(n5131), .A1(n5130), .B0(n5129), .Y(n5134) );
  AOI211XL U3689 ( .A0(n5698), .A1(n5603), .B0(n6123), .C0(n6028), .Y(n5128)
         );
  OAI21XL U3690 ( .A0(n4965), .A1(n5093), .B0(n5092), .Y(n4974) );
  AOI211XL U3691 ( .A0(N2758), .A1(n4964), .B0(n5086), .C0(n4963), .Y(n4965)
         );
  AOI211XL U3692 ( .A0(n4962), .A1(n5084), .B0(n5091), .C0(n5083), .Y(n4963)
         );
  AOI31XL U3693 ( .A0(n6124), .A1(n5098), .A2(n5087), .B0(n5085), .Y(n4962) );
  AOI31XL U3694 ( .A0(n6123), .A1(n5098), .A2(n5110), .B0(n5109), .Y(n4875) );
  AOI22XL U3695 ( .A0(N2773), .A1(n4981), .B0(N2774), .B1(n4785), .Y(n5117) );
  AOI21XL U3696 ( .A0(N2781), .A1(n4971), .B0(N2782), .Y(n4785) );
  AOI2BB2XL U3697 ( .B0(n5698), .B1(n4985), .A0N(n4872), .A1N(n8569), .Y(n5154) );
  OAI22XL U3698 ( .A0(N2766), .A1(n5704), .B0(n8568), .B1(n4979), .Y(n5156) );
  AOI22XL U3699 ( .A0(N2766), .A1(n5704), .B0(N2765), .B1(n4981), .Y(n5155) );
  AOI2BB2XL U3700 ( .B0(N2781), .B1(n4989), .A0N(n5807), .A1N(n8567), .Y(n5159) );
  AOI22XL U3701 ( .A0(n6123), .A1(n6028), .B0(n5698), .B1(n5603), .Y(n4980) );
  OAI22XL U3702 ( .A0(N2758), .A1(n5704), .B0(N2757), .B1(n4981), .Y(n5129) );
  CLKINVX3 U3703 ( .A(n3450), .Y(n4959) );
  CLKINVX3 U3704 ( .A(n5165), .Y(n4777) );
  AOI22XL U3705 ( .A0(n6498), .A1(n6073), .B0(n6072), .B1(n6495), .Y(n6120) );
  AOI22XL U3706 ( .A0(n6574), .A1(n6115), .B0(n6114), .B1(n6571), .Y(n6119) );
  NOR4XL U3707 ( .A(n6051), .B(n6050), .C(n6049), .D(n6048), .Y(n6073) );
  AOI22XL U3708 ( .A0(n6498), .A1(n5649), .B0(n5648), .B1(n6495), .Y(n5695) );
  AOI22XL U3709 ( .A0(n6574), .A1(n5691), .B0(n5690), .B1(n6571), .Y(n5694) );
  NOR4XL U3710 ( .A(n5627), .B(n5626), .C(n5625), .D(n5624), .Y(n5649) );
  AOI22XL U3711 ( .A0(n6498), .A1(n6497), .B0(n6496), .B1(n6495), .Y(n6580) );
  NOR4XL U3712 ( .A(n6442), .B(n6441), .C(n6440), .D(n6439), .Y(n6497) );
  NOR4XL U3713 ( .A(n6494), .B(n6493), .C(n6492), .D(n6491), .Y(n6496) );
  NAND4XL U3714 ( .A(n6438), .B(n6437), .C(n6436), .D(n6435), .Y(n6439) );
  AOI31XL U3715 ( .A0(n6127), .A1(n5084), .A2(n6028), .B0(n5083), .Y(n5088) );
  NAND2XL U3716 ( .A(n4871), .B(n5603), .Y(n5087) );
  NOR2XL U3717 ( .A(N2776), .B(n4986), .Y(n5085) );
  NOR2XL U3718 ( .A(N2775), .B(n6173), .Y(n5086) );
  NOR2XL U3719 ( .A(N2759), .B(n4967), .Y(n5091) );
  AOI31XL U3720 ( .A0(n6126), .A1(n5098), .A2(n5097), .B0(n5099), .Y(n4969) );
  AOI22XL U3721 ( .A0(n8569), .A1(n4872), .B0(n8568), .B1(n4979), .Y(n5151) );
  INVXL U3722 ( .A(N2784), .Y(n4872) );
  INVX1 U3723 ( .A(n5194), .Y(n5192) );
  INVXL U3724 ( .A(n5214), .Y(n5208) );
  AOI22XL U3725 ( .A0(n5117), .A1(n5116), .B0(N2780), .B1(n5115), .Y(n5121) );
  AOI21XL U3726 ( .A0(n5111), .A1(n5110), .B0(n5109), .Y(n5114) );
  NAND2XL U3727 ( .A(n6127), .B(n6029), .Y(n5111) );
  AOI21XL U3728 ( .A0(n5105), .A1(n5104), .B0(n5103), .Y(n5108) );
  OAI31XL U3729 ( .A0(n5099), .A1(n6126), .A2(n5098), .B0(n5097), .Y(n5101) );
  OAI22XL U3730 ( .A0(n8567), .A1(n5115), .B0(N2765), .B1(n4971), .Y(n5107) );
  INVXL U3731 ( .A(n5151), .Y(n5152) );
  OAI31XL U3732 ( .A0(n6126), .A1(n5136), .A2(n6028), .B0(n5135), .Y(n5138) );
  AOI22XL U3733 ( .A0(n6401), .A1(n5011), .B0(n5014), .B1(n8524), .Y(n5006) );
  INVXL U3734 ( .A(n5042), .Y(n5036) );
  OAI22XL U3735 ( .A0(N2779), .A1(n5118), .B0(N2780), .B1(n5115), .Y(n5120) );
  OAI21XL U3736 ( .A0(n4972), .A1(n5107), .B0(n5106), .Y(n4973) );
  AOI21XL U3737 ( .A0(n5105), .A1(n4970), .B0(n5103), .Y(n4972) );
  AOI22XL U3738 ( .A0(n4969), .A1(n5100), .B0(n5102), .B1(n4968), .Y(n4970) );
  NAND2XL U3739 ( .A(n8568), .B(n4967), .Y(n4968) );
  AOI22XL U3740 ( .A0(N2771), .A1(n4993), .B0(N2772), .B1(n5806), .Y(n5096) );
  INVX1 U3741 ( .A(N2771), .Y(n5118) );
  NAND2XL U3742 ( .A(N2771), .B(n3441), .Y(n5124) );
  AOI22XL U3743 ( .A0(N2758), .A1(n5704), .B0(N2759), .B1(n4979), .Y(n5131) );
  AOI22XL U3744 ( .A0(n4988), .A1(n5137), .B0(n5139), .B1(n4987), .Y(n4991) );
  NAND2XL U3745 ( .A(n8568), .B(n6173), .Y(n4987) );
  AOI31XL U3746 ( .A0(n6126), .A1(n6028), .A2(n5135), .B0(n5136), .Y(n4988) );
  AOI22XL U3747 ( .A0(n8567), .A1(n5806), .B0(n3442), .B1(n4993), .Y(n5143) );
  OAI22XL U3748 ( .A0(n8567), .A1(n5806), .B0(N2765), .B1(n4992), .Y(n5144) );
  OAI22XL U3749 ( .A0(N2780), .A1(n5806), .B0(N2781), .B1(n4992), .Y(n5133) );
  AOI22XL U3750 ( .A0(N2780), .A1(n5806), .B0(N2779), .B1(n4993), .Y(n5132) );
  OAI21XL U3751 ( .A0(n5162), .A1(n4784), .B0(n5160), .Y(n4997) );
  AOI22XL U3752 ( .A0(n5159), .A1(n4783), .B0(n8567), .B1(n5807), .Y(n4784) );
  AOI31XL U3753 ( .A0(n6126), .A1(n5154), .A2(n6029), .B0(n4781), .Y(n4782) );
  INVX1 U3754 ( .A(n5177), .Y(n5185) );
  INVX1 U3755 ( .A(n5179), .Y(n5182) );
  NOR2BXL U3756 ( .AN(n5164), .B(n5163), .Y(n5183) );
  NOR2BXL U3757 ( .AN(n5166), .B(n5185), .Y(n5187) );
  AOI22XL U3758 ( .A0(n3935), .A1(image_data[371]), .B0(n3799), .B1(
        image_data[499]), .Y(n3733) );
  AOI22XL U3759 ( .A0(n3798), .A1(image_data[307]), .B0(n3936), .B1(
        image_data[435]), .Y(n3734) );
  AOI22XL U3760 ( .A0(n3884), .A1(image_data[275]), .B0(n3934), .B1(
        image_data[403]), .Y(n3736) );
  AOI22XL U3761 ( .A0(n3885), .A1(image_data[339]), .B0(n3797), .B1(
        image_data[467]), .Y(n3735) );
  NAND4XL U3762 ( .A(n3764), .B(n3763), .C(n3762), .D(n3761), .Y(n3765) );
  AOI22XL U3763 ( .A0(n3875), .A1(image_data[91]), .B0(n3810), .B1(
        image_data[219]), .Y(n3763) );
  AOI22XL U3764 ( .A0(n3877), .A1(image_data[59]), .B0(n3949), .B1(
        image_data[187]), .Y(n3762) );
  AOI22XL U3765 ( .A0(n3874), .A1(image_data[27]), .B0(n3948), .B1(
        image_data[155]), .Y(n3764) );
  NAND4XL U3766 ( .A(n3752), .B(n3751), .C(n3750), .D(n3749), .Y(n3768) );
  AOI22XL U3767 ( .A0(n3791), .A1(image_data[35]), .B0(n3929), .B1(
        image_data[163]), .Y(n3750) );
  AOI22XL U3768 ( .A0(n3897), .A1(image_data[3]), .B0(n3896), .B1(
        image_data[131]), .Y(n3752) );
  AOI22XL U3769 ( .A0(n3895), .A1(image_data[67]), .B0(n3364), .B1(
        image_data[195]), .Y(n3751) );
  NAND4XL U3770 ( .A(n3760), .B(n3759), .C(n3758), .D(n3757), .Y(n3766) );
  AOI22XL U3771 ( .A0(n3866), .A1(image_data[75]), .B0(n3804), .B1(
        image_data[203]), .Y(n3759) );
  AOI22XL U3772 ( .A0(n3865), .A1(image_data[11]), .B0(n3941), .B1(
        image_data[139]), .Y(n3760) );
  AOI22XL U3773 ( .A0(n3942), .A1(image_data[43]), .B0(n3943), .B1(
        image_data[171]), .Y(n3758) );
  NAND4XL U3774 ( .A(n3756), .B(n3755), .C(n3754), .D(n3753), .Y(n3767) );
  AOI22XL U3775 ( .A0(n3885), .A1(image_data[83]), .B0(n3797), .B1(
        image_data[211]), .Y(n3755) );
  AOI22XL U3776 ( .A0(n3884), .A1(image_data[19]), .B0(n3934), .B1(
        image_data[147]), .Y(n3756) );
  AOI22XL U3777 ( .A0(n3798), .A1(image_data[51]), .B0(n3936), .B1(
        image_data[179]), .Y(n3754) );
  NAND4XL U3778 ( .A(n3744), .B(n3743), .C(n3742), .D(n3741), .Y(n3745) );
  AOI22XL U3779 ( .A0(n3875), .A1(image_data[347]), .B0(n3810), .B1(
        image_data[475]), .Y(n3743) );
  AOI22XL U3780 ( .A0(n3877), .A1(image_data[315]), .B0(n3949), .B1(
        image_data[443]), .Y(n3742) );
  AOI22XL U3781 ( .A0(n3874), .A1(image_data[283]), .B0(n3948), .B1(
        image_data[411]), .Y(n3744) );
  NAND4XL U3782 ( .A(n3732), .B(n3731), .C(n3730), .D(n3729), .Y(n3748) );
  AOI22XL U3783 ( .A0(n3791), .A1(image_data[291]), .B0(n3929), .B1(
        image_data[419]), .Y(n3730) );
  AOI22XL U3784 ( .A0(n3897), .A1(image_data[259]), .B0(n3896), .B1(
        image_data[387]), .Y(n3732) );
  AOI22XL U3785 ( .A0(n3895), .A1(image_data[323]), .B0(n3364), .B1(
        image_data[451]), .Y(n3731) );
  NAND4XL U3786 ( .A(n3740), .B(n3739), .C(n3738), .D(n3737), .Y(n3746) );
  AOI22XL U3787 ( .A0(n3866), .A1(image_data[331]), .B0(n3804), .B1(
        image_data[459]), .Y(n3739) );
  AOI22XL U3788 ( .A0(n3865), .A1(image_data[267]), .B0(n3941), .B1(
        image_data[395]), .Y(n3740) );
  AOI22XL U3789 ( .A0(n3942), .A1(image_data[299]), .B0(n3943), .B1(
        image_data[427]), .Y(n3738) );
  NAND4XL U3790 ( .A(n3511), .B(n3510), .C(n3509), .D(n3508), .Y(n3512) );
  AOI22XL U3791 ( .A0(n3876), .A1(image_data[31]), .B0(n3875), .B1(
        image_data[159]), .Y(n3511) );
  AOI22XL U3792 ( .A0(n3879), .A1(image_data[63]), .B0(n3878), .B1(
        image_data[191]), .Y(n3509) );
  AOI22XL U3793 ( .A0(n3877), .A1(image_data[127]), .B0(n3949), .B1(
        image_data[255]), .Y(n3508) );
  NAND4XL U3794 ( .A(n3507), .B(n3506), .C(n3505), .D(n3504), .Y(n3513) );
  AOI22XL U3795 ( .A0(n3867), .A1(image_data[15]), .B0(n3866), .B1(
        image_data[143]), .Y(n3507) );
  AOI22XL U3796 ( .A0(n3865), .A1(image_data[79]), .B0(n3941), .B1(
        image_data[207]), .Y(n3506) );
  AOI22XL U3797 ( .A0(n3869), .A1(image_data[47]), .B0(n3868), .B1(
        image_data[175]), .Y(n3505) );
  NAND4XL U3798 ( .A(n3503), .B(n3502), .C(n3501), .D(n3500), .Y(n3514) );
  AOI22XL U3799 ( .A0(n3888), .A1(image_data[55]), .B0(n4763), .B1(
        image_data[183]), .Y(n3501) );
  AOI22XL U3800 ( .A0(n3886), .A1(image_data[23]), .B0(n3885), .B1(
        image_data[151]), .Y(n3503) );
  AOI22XL U3801 ( .A0(n3887), .A1(image_data[119]), .B0(n3936), .B1(
        image_data[247]), .Y(n3500) );
  NAND4XL U3802 ( .A(n3499), .B(n3498), .C(n3497), .D(n3496), .Y(n3515) );
  AOI22XL U3803 ( .A0(n3364), .A1(image_data[7]), .B0(n4681), .B1(
        image_data[135]), .Y(n3499) );
  AOI22XL U3804 ( .A0(n3897), .A1(image_data[71]), .B0(n3896), .B1(
        image_data[199]), .Y(n3498) );
  AOI22XL U3805 ( .A0(n3928), .A1(image_data[103]), .B0(n3929), .B1(
        image_data[231]), .Y(n3496) );
  NAND4XL U3806 ( .A(n3491), .B(n3490), .C(n3489), .D(n3488), .Y(n3492) );
  AOI22XL U3807 ( .A0(n3876), .A1(image_data[287]), .B0(n3875), .B1(
        image_data[415]), .Y(n3491) );
  AOI22XL U3808 ( .A0(n3879), .A1(image_data[319]), .B0(n3878), .B1(
        image_data[447]), .Y(n3489) );
  AOI22XL U3809 ( .A0(n3877), .A1(image_data[383]), .B0(n3949), .B1(
        image_data[511]), .Y(n3488) );
  NAND4XL U3810 ( .A(n3480), .B(n3479), .C(n3478), .D(n3477), .Y(n3493) );
  AOI22XL U3811 ( .A0(n3867), .A1(image_data[271]), .B0(n3866), .B1(
        image_data[399]), .Y(n3480) );
  AOI22XL U3812 ( .A0(n4753), .A1(image_data[335]), .B0(n3941), .B1(
        image_data[463]), .Y(n3479) );
  AOI22XL U3813 ( .A0(n3869), .A1(image_data[303]), .B0(n3868), .B1(
        image_data[431]), .Y(n3478) );
  NAND4XL U3814 ( .A(n3475), .B(n3474), .C(n3473), .D(n3472), .Y(n3494) );
  AOI22XL U3815 ( .A0(n3888), .A1(image_data[311]), .B0(n4763), .B1(
        image_data[439]), .Y(n3473) );
  AOI22XL U3816 ( .A0(n3886), .A1(image_data[279]), .B0(n3885), .B1(
        image_data[407]), .Y(n3475) );
  AOI22XL U3817 ( .A0(n3887), .A1(image_data[375]), .B0(n3936), .B1(
        image_data[503]), .Y(n3472) );
  NAND4XL U3818 ( .A(n3469), .B(n3468), .C(n3467), .D(n3466), .Y(n3495) );
  AOI22XL U3819 ( .A0(n3364), .A1(image_data[263]), .B0(n4681), .B1(
        image_data[391]), .Y(n3469) );
  AOI22XL U3820 ( .A0(n3897), .A1(image_data[327]), .B0(n3896), .B1(
        image_data[455]), .Y(n3468) );
  AOI22XL U3821 ( .A0(n3928), .A1(image_data[359]), .B0(n3929), .B1(
        image_data[487]), .Y(n3466) );
  INVX1 U3822 ( .A(n5007), .Y(n5015) );
  AND2X1 U3823 ( .A(n4998), .B(n4997), .Y(n5011) );
  NOR2BXL U3824 ( .AN(n4999), .B(n5015), .Y(n5014) );
  AOI22XL U3825 ( .A0(n3879), .A1(image_data[306]), .B0(n3878), .B1(
        image_data[434]), .Y(n3827) );
  AOI22XL U3826 ( .A0(n3874), .A1(image_data[338]), .B0(n3948), .B1(
        image_data[466]), .Y(n3828) );
  AOI22XL U3827 ( .A0(n3877), .A1(image_data[370]), .B0(n3949), .B1(
        image_data[498]), .Y(n3826) );
  AOI22XL U3828 ( .A0(n3876), .A1(image_data[274]), .B0(n3875), .B1(
        image_data[402]), .Y(n3829) );
  NAND4XL U3829 ( .A(n3857), .B(n3856), .C(n3855), .D(n3854), .Y(n3858) );
  AOI22XL U3830 ( .A0(n3928), .A1(image_data[90]), .B0(n3929), .B1(
        image_data[218]), .Y(n3856) );
  AOI22XL U3831 ( .A0(n3897), .A1(image_data[58]), .B0(n3896), .B1(
        image_data[186]), .Y(n3855) );
  AOI22XL U3832 ( .A0(n3894), .A1(image_data[26]), .B0(n3893), .B1(
        image_data[154]), .Y(n3857) );
  NAND4XL U3833 ( .A(n3853), .B(n3852), .C(n3851), .D(n3850), .Y(n3859) );
  AOI22XL U3834 ( .A0(n3886), .A1(image_data[10]), .B0(n3885), .B1(
        image_data[138]), .Y(n3853) );
  AOI22XL U3835 ( .A0(n3887), .A1(image_data[106]), .B0(n3936), .B1(
        image_data[234]), .Y(n3850) );
  AOI22XL U3836 ( .A0(n3884), .A1(image_data[74]), .B0(n3934), .B1(
        image_data[202]), .Y(n3852) );
  NAND4XL U3837 ( .A(n3845), .B(n3844), .C(n3843), .D(n3842), .Y(n3861) );
  AOI22XL U3838 ( .A0(n3865), .A1(image_data[66]), .B0(n3941), .B1(
        image_data[194]), .Y(n3844) );
  AOI22XL U3839 ( .A0(n3867), .A1(image_data[2]), .B0(n3866), .B1(
        image_data[130]), .Y(n3845) );
  AOI22XL U3840 ( .A0(n3942), .A1(image_data[98]), .B0(n3943), .B1(
        image_data[226]), .Y(n3842) );
  NAND4XL U3841 ( .A(n3849), .B(n3848), .C(n3847), .D(n3846), .Y(n3860) );
  AOI22XL U3842 ( .A0(n3876), .A1(image_data[18]), .B0(n3875), .B1(
        image_data[146]), .Y(n3849) );
  AOI22XL U3843 ( .A0(n3877), .A1(image_data[114]), .B0(n3949), .B1(
        image_data[242]), .Y(n3846) );
  AOI22XL U3844 ( .A0(n3874), .A1(image_data[82]), .B0(n3948), .B1(
        image_data[210]), .Y(n3848) );
  NAND4XL U3845 ( .A(n3837), .B(n3836), .C(n3835), .D(n3834), .Y(n3838) );
  AOI22XL U3846 ( .A0(n4670), .A1(image_data[314]), .B0(n3896), .B1(
        image_data[442]), .Y(n3835) );
  AOI22XL U3847 ( .A0(n3928), .A1(image_data[346]), .B0(n3929), .B1(
        image_data[474]), .Y(n3836) );
  AOI22XL U3848 ( .A0(n3894), .A1(image_data[282]), .B0(n3893), .B1(
        image_data[410]), .Y(n3837) );
  NAND4XL U3849 ( .A(n3833), .B(n3832), .C(n3831), .D(n3830), .Y(n3839) );
  AOI22XL U3850 ( .A0(n3886), .A1(image_data[266]), .B0(n3885), .B1(
        image_data[394]), .Y(n3833) );
  AOI22XL U3851 ( .A0(n3887), .A1(image_data[362]), .B0(n3936), .B1(
        image_data[490]), .Y(n3830) );
  AOI22XL U3852 ( .A0(n3884), .A1(image_data[330]), .B0(n3934), .B1(
        image_data[458]), .Y(n3832) );
  NAND4XL U3853 ( .A(n3825), .B(n3824), .C(n3823), .D(n3822), .Y(n3841) );
  AOI22XL U3854 ( .A0(n3865), .A1(image_data[322]), .B0(n3941), .B1(
        image_data[450]), .Y(n3824) );
  AOI22XL U3855 ( .A0(n3867), .A1(image_data[258]), .B0(n3866), .B1(
        image_data[386]), .Y(n3825) );
  AOI22XL U3856 ( .A0(n3942), .A1(image_data[354]), .B0(n3943), .B1(
        image_data[482]), .Y(n3822) );
  AOI22XL U3857 ( .A0(n3935), .A1(image_data[372]), .B0(n3888), .B1(
        image_data[500]), .Y(n4455) );
  AOI22XL U3858 ( .A0(n3887), .A1(image_data[308]), .B0(n3936), .B1(
        image_data[436]), .Y(n4456) );
  NAND4XL U3859 ( .A(n4486), .B(n4485), .C(n4484), .D(n4483), .Y(n4487) );
  AOI22XL U3860 ( .A0(n3875), .A1(image_data[92]), .B0(n3876), .B1(
        image_data[220]), .Y(n4485) );
  AOI22XL U3861 ( .A0(n3877), .A1(image_data[60]), .B0(n3949), .B1(
        image_data[188]), .Y(n4484) );
  AOI22XL U3862 ( .A0(n3874), .A1(image_data[28]), .B0(n3948), .B1(
        image_data[156]), .Y(n4486) );
  NAND4XL U3863 ( .A(n4482), .B(n4481), .C(n4480), .D(n4479), .Y(n4488) );
  AOI22XL U3864 ( .A0(n3866), .A1(image_data[76]), .B0(n3867), .B1(
        image_data[204]), .Y(n4481) );
  AOI22XL U3865 ( .A0(n3865), .A1(image_data[12]), .B0(n3941), .B1(
        image_data[140]), .Y(n4482) );
  AOI22XL U3866 ( .A0(n3942), .A1(image_data[44]), .B0(n3943), .B1(
        image_data[172]), .Y(n4480) );
  NAND4XL U3867 ( .A(n4474), .B(n4473), .C(n4472), .D(n4471), .Y(n4490) );
  AOI22XL U3868 ( .A0(n3897), .A1(image_data[4]), .B0(n3896), .B1(
        image_data[132]), .Y(n4474) );
  AOI22XL U3869 ( .A0(n3928), .A1(image_data[36]), .B0(n3929), .B1(
        image_data[164]), .Y(n4472) );
  AOI22XL U3870 ( .A0(n3895), .A1(image_data[68]), .B0(n3364), .B1(
        image_data[196]), .Y(n4473) );
  NAND4XL U3871 ( .A(n4478), .B(n4477), .C(n4476), .D(n4475), .Y(n4489) );
  AOI22XL U3872 ( .A0(n3885), .A1(image_data[84]), .B0(n3886), .B1(
        image_data[212]), .Y(n4477) );
  AOI22XL U3873 ( .A0(n3884), .A1(image_data[20]), .B0(n3934), .B1(
        image_data[148]), .Y(n4478) );
  AOI22XL U3874 ( .A0(n3887), .A1(image_data[52]), .B0(n3936), .B1(
        image_data[180]), .Y(n4476) );
  NAND4XL U3875 ( .A(n4466), .B(n4465), .C(n4464), .D(n4463), .Y(n4467) );
  AOI22XL U3876 ( .A0(n3875), .A1(image_data[348]), .B0(n3876), .B1(
        image_data[476]), .Y(n4465) );
  AOI22XL U3877 ( .A0(n3877), .A1(image_data[316]), .B0(n3949), .B1(
        image_data[444]), .Y(n4464) );
  AOI22XL U3878 ( .A0(n3874), .A1(image_data[284]), .B0(n3948), .B1(
        image_data[412]), .Y(n4466) );
  NAND4XL U3879 ( .A(n4462), .B(n4461), .C(n4460), .D(n4459), .Y(n4468) );
  AOI22XL U3880 ( .A0(n3865), .A1(image_data[268]), .B0(n3941), .B1(
        image_data[396]), .Y(n4462) );
  AOI22XL U3881 ( .A0(n3866), .A1(image_data[332]), .B0(n3867), .B1(
        image_data[460]), .Y(n4461) );
  AOI22XL U3882 ( .A0(n3942), .A1(image_data[300]), .B0(n3943), .B1(
        image_data[428]), .Y(n4460) );
  NAND4XL U3883 ( .A(n4454), .B(n4453), .C(n4452), .D(n4451), .Y(n4470) );
  AOI22XL U3884 ( .A0(n3897), .A1(image_data[260]), .B0(n3896), .B1(
        image_data[388]), .Y(n4454) );
  AOI22XL U3885 ( .A0(n3928), .A1(image_data[292]), .B0(n3929), .B1(
        image_data[420]), .Y(n4452) );
  AOI22XL U3886 ( .A0(n3895), .A1(image_data[324]), .B0(n3364), .B1(
        image_data[452]), .Y(n4453) );
  AOI22XL U3887 ( .A0(n3894), .A1(image_data[284]), .B0(n3893), .B1(
        image_data[412]), .Y(n3659) );
  AOI22XL U3888 ( .A0(n3928), .A1(image_data[348]), .B0(n3929), .B1(
        image_data[476]), .Y(n3658) );
  AOI22XL U3889 ( .A0(n3897), .A1(image_data[316]), .B0(n3896), .B1(
        image_data[444]), .Y(n3657) );
  AOI22XL U3890 ( .A0(n4681), .A1(image_data[380]), .B0(n3364), .B1(
        image_data[508]), .Y(n3656) );
  NAND4XL U3891 ( .A(n3679), .B(n3678), .C(n3677), .D(n3676), .Y(n3680) );
  AOI22XL U3892 ( .A0(n3897), .A1(image_data[60]), .B0(n3896), .B1(
        image_data[188]), .Y(n3677) );
  AOI22XL U3893 ( .A0(n3928), .A1(image_data[92]), .B0(n3929), .B1(
        image_data[220]), .Y(n3678) );
  AOI22XL U3894 ( .A0(n3894), .A1(image_data[28]), .B0(n3893), .B1(
        image_data[156]), .Y(n3679) );
  NAND4XL U3895 ( .A(n3675), .B(n3674), .C(n3673), .D(n3672), .Y(n3681) );
  AOI22XL U3896 ( .A0(n3886), .A1(image_data[12]), .B0(n3885), .B1(
        image_data[140]), .Y(n3675) );
  AOI22XL U3897 ( .A0(n3887), .A1(image_data[108]), .B0(n3936), .B1(
        image_data[236]), .Y(n3672) );
  AOI22XL U3898 ( .A0(n3884), .A1(image_data[76]), .B0(n3934), .B1(
        image_data[204]), .Y(n3674) );
  NAND4XL U3899 ( .A(n3667), .B(n3666), .C(n3665), .D(n3664), .Y(n3683) );
  AOI22XL U3900 ( .A0(n3867), .A1(image_data[4]), .B0(n3866), .B1(
        image_data[132]), .Y(n3667) );
  AOI22XL U3901 ( .A0(n3865), .A1(image_data[68]), .B0(n3941), .B1(
        image_data[196]), .Y(n3666) );
  AOI22XL U3902 ( .A0(n3942), .A1(image_data[100]), .B0(n3943), .B1(
        image_data[228]), .Y(n3664) );
  NAND4XL U3903 ( .A(n3671), .B(n3670), .C(n3669), .D(n3668), .Y(n3682) );
  AOI22XL U3904 ( .A0(n3876), .A1(image_data[20]), .B0(n3875), .B1(
        image_data[148]), .Y(n3671) );
  AOI22XL U3905 ( .A0(n3877), .A1(image_data[116]), .B0(n3949), .B1(
        image_data[244]), .Y(n3668) );
  AOI22XL U3906 ( .A0(n3874), .A1(image_data[84]), .B0(n3948), .B1(
        image_data[212]), .Y(n3670) );
  NAND4XL U3907 ( .A(n3655), .B(n3654), .C(n3653), .D(n3652), .Y(n3661) );
  AOI22XL U3908 ( .A0(n3886), .A1(image_data[268]), .B0(n3885), .B1(
        image_data[396]), .Y(n3655) );
  AOI22XL U3909 ( .A0(n3887), .A1(image_data[364]), .B0(n3936), .B1(
        image_data[492]), .Y(n3652) );
  AOI22XL U3910 ( .A0(n3884), .A1(image_data[332]), .B0(n3934), .B1(
        image_data[460]), .Y(n3654) );
  NAND4XL U3911 ( .A(n3647), .B(n3646), .C(n3645), .D(n3644), .Y(n3663) );
  AOI22XL U3912 ( .A0(n3867), .A1(image_data[260]), .B0(n3866), .B1(
        image_data[388]), .Y(n3647) );
  AOI22XL U3913 ( .A0(n3865), .A1(image_data[324]), .B0(n3941), .B1(
        image_data[452]), .Y(n3646) );
  AOI22XL U3914 ( .A0(n3942), .A1(image_data[356]), .B0(n3943), .B1(
        image_data[484]), .Y(n3644) );
  NAND4XL U3915 ( .A(n3651), .B(n3650), .C(n3649), .D(n3648), .Y(n3662) );
  AOI22XL U3916 ( .A0(n3876), .A1(image_data[276]), .B0(n3875), .B1(
        image_data[404]), .Y(n3651) );
  AOI22XL U3917 ( .A0(n3877), .A1(image_data[372]), .B0(n3949), .B1(
        image_data[500]), .Y(n3648) );
  AOI22XL U3918 ( .A0(n3874), .A1(image_data[340]), .B0(n3948), .B1(
        image_data[468]), .Y(n3650) );
  AOI22XL U3919 ( .A0(n4721), .A1(image_data[371]), .B0(n3879), .B1(
        image_data[499]), .Y(n4280) );
  AOI22XL U3920 ( .A0(n3874), .A1(image_data[275]), .B0(n3948), .B1(
        image_data[403]), .Y(n4283) );
  AOI22XL U3921 ( .A0(n3877), .A1(image_data[307]), .B0(n3949), .B1(
        image_data[435]), .Y(n4281) );
  AOI22XL U3922 ( .A0(n4719), .A1(image_data[339]), .B0(n3876), .B1(
        image_data[467]), .Y(n4282) );
  NAND4XL U3923 ( .A(n4311), .B(n4310), .C(n4309), .D(n4308), .Y(n4312) );
  AOI22XL U3924 ( .A0(n3928), .A1(image_data[27]), .B0(n3929), .B1(
        image_data[155]), .Y(n4311) );
  AOI22XL U3925 ( .A0(n3896), .A1(image_data[123]), .B0(n3897), .B1(
        image_data[251]), .Y(n4308) );
  AOI22XL U3926 ( .A0(n4702), .A1(image_data[91]), .B0(n3894), .B1(
        image_data[219]), .Y(n4310) );
  NAND4XL U3927 ( .A(n4307), .B(n4306), .C(n4305), .D(n4304), .Y(n4313) );
  AOI22XL U3928 ( .A0(n4707), .A1(image_data[75]), .B0(n3886), .B1(
        image_data[203]), .Y(n4306) );
  AOI22XL U3929 ( .A0(n3884), .A1(image_data[11]), .B0(n3934), .B1(
        image_data[139]), .Y(n4307) );
  AOI22XL U3930 ( .A0(n3887), .A1(image_data[43]), .B0(n3936), .B1(
        image_data[171]), .Y(n4305) );
  NAND4XL U3931 ( .A(n4303), .B(n4302), .C(n4301), .D(n4300), .Y(n4314) );
  AOI22XL U3932 ( .A0(n4719), .A1(image_data[83]), .B0(n3876), .B1(
        image_data[211]), .Y(n4302) );
  AOI22XL U3933 ( .A0(n3877), .A1(image_data[51]), .B0(n3949), .B1(
        image_data[179]), .Y(n4301) );
  AOI22XL U3934 ( .A0(n3874), .A1(image_data[19]), .B0(n3948), .B1(
        image_data[147]), .Y(n4303) );
  NAND4XL U3935 ( .A(n4299), .B(n4298), .C(n4297), .D(n4296), .Y(n4315) );
  AOI22XL U3936 ( .A0(n3865), .A1(image_data[3]), .B0(n3941), .B1(
        image_data[131]), .Y(n4299) );
  AOI22XL U3937 ( .A0(n3866), .A1(image_data[67]), .B0(n3867), .B1(
        image_data[195]), .Y(n4298) );
  AOI22XL U3938 ( .A0(n3942), .A1(image_data[35]), .B0(n3943), .B1(
        image_data[163]), .Y(n4297) );
  NAND4XL U3939 ( .A(n4291), .B(n4290), .C(n4289), .D(n4288), .Y(n4292) );
  AOI22XL U3940 ( .A0(n3928), .A1(image_data[283]), .B0(n3929), .B1(
        image_data[411]), .Y(n4291) );
  AOI22XL U3941 ( .A0(n3896), .A1(image_data[379]), .B0(n3897), .B1(
        image_data[507]), .Y(n4288) );
  AOI22XL U3942 ( .A0(n4702), .A1(image_data[347]), .B0(n3894), .B1(
        image_data[475]), .Y(n4290) );
  NAND4XL U3943 ( .A(n4279), .B(n4278), .C(n4277), .D(n4276), .Y(n4295) );
  AOI22XL U3944 ( .A0(n3865), .A1(image_data[259]), .B0(n3941), .B1(
        image_data[387]), .Y(n4279) );
  AOI22XL U3945 ( .A0(n3866), .A1(image_data[323]), .B0(n3867), .B1(
        image_data[451]), .Y(n4278) );
  AOI22XL U3946 ( .A0(n3942), .A1(image_data[291]), .B0(n3943), .B1(
        image_data[419]), .Y(n4277) );
  NAND4XL U3947 ( .A(n4287), .B(n4286), .C(n4285), .D(n4284), .Y(n4293) );
  AOI22XL U3948 ( .A0(n4707), .A1(image_data[331]), .B0(n3886), .B1(
        image_data[459]), .Y(n4286) );
  AOI22XL U3949 ( .A0(n3884), .A1(image_data[267]), .B0(n3934), .B1(
        image_data[395]), .Y(n4287) );
  AOI22XL U3950 ( .A0(n3887), .A1(image_data[299]), .B0(n3936), .B1(
        image_data[427]), .Y(n4285) );
  AOI22XL U3951 ( .A0(n3942), .A1(image_data[288]), .B0(n3943), .B1(
        image_data[416]), .Y(n4787) );
  AOI22XL U3952 ( .A0(n4714), .A1(image_data[352]), .B0(n3869), .B1(
        image_data[480]), .Y(n4786) );
  AOI22XL U3953 ( .A0(n3865), .A1(image_data[256]), .B0(n3941), .B1(
        image_data[384]), .Y(n4789) );
  AOI22XL U3954 ( .A0(n3866), .A1(image_data[320]), .B0(n3867), .B1(
        image_data[448]), .Y(n4788) );
  NAND4XL U3955 ( .A(n4821), .B(n4820), .C(n4819), .D(n4818), .Y(n4822) );
  AOI22XL U3956 ( .A0(n4702), .A1(image_data[88]), .B0(n3894), .B1(
        image_data[216]), .Y(n4820) );
  AOI22XL U3957 ( .A0(n3896), .A1(image_data[120]), .B0(n3897), .B1(
        image_data[248]), .Y(n4818) );
  AOI22XL U3958 ( .A0(n3928), .A1(image_data[24]), .B0(n3929), .B1(
        image_data[152]), .Y(n4821) );
  NAND4XL U3959 ( .A(n4817), .B(n4816), .C(n4815), .D(n4814), .Y(n4823) );
  AOI22XL U3960 ( .A0(n3885), .A1(image_data[72]), .B0(n3886), .B1(
        image_data[200]), .Y(n4816) );
  AOI22XL U3961 ( .A0(n3884), .A1(image_data[8]), .B0(n3934), .B1(
        image_data[136]), .Y(n4817) );
  AOI22XL U3962 ( .A0(n3887), .A1(image_data[40]), .B0(n3936), .B1(
        image_data[168]), .Y(n4815) );
  NAND4XL U3963 ( .A(n4813), .B(n4812), .C(n4811), .D(n4810), .Y(n4824) );
  AOI22XL U3964 ( .A0(n4719), .A1(image_data[80]), .B0(n3876), .B1(
        image_data[208]), .Y(n4812) );
  AOI22XL U3965 ( .A0(n4721), .A1(image_data[112]), .B0(n3879), .B1(
        image_data[240]), .Y(n4810) );
  AOI22XL U3966 ( .A0(n3877), .A1(image_data[48]), .B0(n3949), .B1(
        image_data[176]), .Y(n4811) );
  NAND4XL U3967 ( .A(n4809), .B(n4808), .C(n4807), .D(n4806), .Y(n4825) );
  AOI22XL U3968 ( .A0(n3866), .A1(image_data[64]), .B0(n3867), .B1(
        image_data[192]), .Y(n4808) );
  AOI22XL U3969 ( .A0(n3865), .A1(image_data[0]), .B0(n3941), .B1(
        image_data[128]), .Y(n4809) );
  AOI22XL U3970 ( .A0(n4714), .A1(image_data[96]), .B0(n3869), .B1(
        image_data[224]), .Y(n4806) );
  NAND4XL U3971 ( .A(n4801), .B(n4800), .C(n4799), .D(n4798), .Y(n4802) );
  AOI22XL U3972 ( .A0(n4702), .A1(image_data[344]), .B0(n3894), .B1(
        image_data[472]), .Y(n4800) );
  AOI22XL U3973 ( .A0(n3896), .A1(image_data[376]), .B0(n3897), .B1(
        image_data[504]), .Y(n4798) );
  AOI22XL U3974 ( .A0(n3928), .A1(image_data[280]), .B0(n3929), .B1(
        image_data[408]), .Y(n4801) );
  NAND4XL U3975 ( .A(n4797), .B(n4796), .C(n4795), .D(n4794), .Y(n4803) );
  AOI22XL U3976 ( .A0(n4707), .A1(image_data[328]), .B0(n3886), .B1(
        image_data[456]), .Y(n4796) );
  AOI22XL U3977 ( .A0(n3884), .A1(image_data[264]), .B0(n3934), .B1(
        image_data[392]), .Y(n4797) );
  AOI22XL U3978 ( .A0(n3887), .A1(image_data[296]), .B0(n3936), .B1(
        image_data[424]), .Y(n4795) );
  NAND4XL U3979 ( .A(n4793), .B(n4792), .C(n4791), .D(n4790), .Y(n4804) );
  AOI22XL U3980 ( .A0(n4719), .A1(image_data[336]), .B0(n3876), .B1(
        image_data[464]), .Y(n4792) );
  AOI22XL U3981 ( .A0(n4721), .A1(image_data[368]), .B0(n3879), .B1(
        image_data[496]), .Y(n4790) );
  AOI22XL U3982 ( .A0(n3877), .A1(image_data[304]), .B0(n3949), .B1(
        image_data[432]), .Y(n4791) );
  NAND4XL U3983 ( .A(n4611), .B(n4610), .C(n4609), .D(n4608), .Y(n4612) );
  AOI22XL U3984 ( .A0(n3876), .A1(image_data[280]), .B0(n4719), .B1(
        image_data[408]), .Y(n4611) );
  AOI22XL U3985 ( .A0(n3879), .A1(image_data[312]), .B0(n4721), .B1(
        image_data[440]), .Y(n4609) );
  AOI22XL U3986 ( .A0(n3877), .A1(image_data[376]), .B0(n3949), .B1(
        image_data[504]), .Y(n4608) );
  NAND4XL U3987 ( .A(n4607), .B(n4606), .C(n4605), .D(n4604), .Y(n4613) );
  AOI22XL U3988 ( .A0(n3869), .A1(image_data[296]), .B0(n4714), .B1(
        image_data[424]), .Y(n4605) );
  AOI22XL U3989 ( .A0(n3867), .A1(image_data[264]), .B0(n3866), .B1(
        image_data[392]), .Y(n4607) );
  AOI22XL U3990 ( .A0(n3865), .A1(image_data[328]), .B0(n3941), .B1(
        image_data[456]), .Y(n4606) );
  NAND4XL U3991 ( .A(n4603), .B(n4602), .C(n4601), .D(n4600), .Y(n4614) );
  AOI22XL U3992 ( .A0(n3886), .A1(image_data[272]), .B0(n4707), .B1(
        image_data[400]), .Y(n4603) );
  AOI22XL U3993 ( .A0(n3887), .A1(image_data[368]), .B0(n3936), .B1(
        image_data[496]), .Y(n4600) );
  AOI22XL U3994 ( .A0(n3888), .A1(image_data[304]), .B0(n3935), .B1(
        image_data[432]), .Y(n4601) );
  NAND4XL U3995 ( .A(n4599), .B(n4598), .C(n4597), .D(n4596), .Y(n4615) );
  AOI22XL U3996 ( .A0(n3894), .A1(image_data[288]), .B0(n4702), .B1(
        image_data[416]), .Y(n4597) );
  AOI22XL U3997 ( .A0(n3364), .A1(image_data[256]), .B0(n4681), .B1(
        image_data[384]), .Y(n4599) );
  AOI22XL U3998 ( .A0(n3897), .A1(image_data[320]), .B0(n3896), .B1(
        image_data[448]), .Y(n4598) );
  NOR4XL U3999 ( .A(n4635), .B(n4634), .C(n4633), .D(n4632), .Y(n4636) );
  NAND4XL U4000 ( .A(n4623), .B(n4622), .C(n4621), .D(n4620), .Y(n4634) );
  NAND4XL U4001 ( .A(n4627), .B(n4626), .C(n4625), .D(n4624), .Y(n4633) );
  NAND4XL U4002 ( .A(n4631), .B(n4630), .C(n4629), .D(n4628), .Y(n4632) );
  AOI22XL U4003 ( .A0(n3935), .A1(image_data[365]), .B0(n3888), .B1(
        image_data[493]), .Y(n4200) );
  AOI22XL U4004 ( .A0(n3887), .A1(image_data[301]), .B0(n3936), .B1(
        image_data[429]), .Y(n4201) );
  AOI22XL U4005 ( .A0(n4708), .A1(image_data[269]), .B0(n3934), .B1(
        image_data[397]), .Y(n4203) );
  AOI22XL U4006 ( .A0(n4707), .A1(image_data[333]), .B0(n3886), .B1(
        image_data[461]), .Y(n4202) );
  NAND4XL U4007 ( .A(n4227), .B(n4226), .C(n4225), .D(n4224), .Y(n4228) );
  AOI22XL U4008 ( .A0(n3896), .A1(image_data[125]), .B0(n3897), .B1(
        image_data[253]), .Y(n4224) );
  AOI22XL U4009 ( .A0(n4702), .A1(image_data[93]), .B0(n3894), .B1(
        image_data[221]), .Y(n4226) );
  AOI22XL U4010 ( .A0(n3928), .A1(image_data[29]), .B0(n3929), .B1(
        image_data[157]), .Y(n4227) );
  NAND4XL U4011 ( .A(n4223), .B(n4222), .C(n4221), .D(n4220), .Y(n4229) );
  AOI22XL U4012 ( .A0(n4707), .A1(image_data[77]), .B0(n3886), .B1(
        image_data[205]), .Y(n4222) );
  AOI22XL U4013 ( .A0(n4708), .A1(image_data[13]), .B0(n3934), .B1(
        image_data[141]), .Y(n4223) );
  AOI22XL U4014 ( .A0(n3887), .A1(image_data[45]), .B0(n3936), .B1(
        image_data[173]), .Y(n4221) );
  NAND4XL U4015 ( .A(n4219), .B(n4218), .C(n4217), .D(n4216), .Y(n4230) );
  AOI22XL U4016 ( .A0(n4719), .A1(image_data[85]), .B0(n3876), .B1(
        image_data[213]), .Y(n4218) );
  AOI22XL U4017 ( .A0(n4721), .A1(image_data[117]), .B0(n3879), .B1(
        image_data[245]), .Y(n4216) );
  AOI22XL U4018 ( .A0(n4722), .A1(image_data[53]), .B0(n3949), .B1(
        image_data[181]), .Y(n4217) );
  NAND4XL U4019 ( .A(n4215), .B(n4214), .C(n4213), .D(n4212), .Y(n4231) );
  AOI22XL U4020 ( .A0(n3865), .A1(image_data[5]), .B0(n3941), .B1(
        image_data[133]), .Y(n4215) );
  AOI22XL U4021 ( .A0(n4714), .A1(image_data[101]), .B0(n3869), .B1(
        image_data[229]), .Y(n4212) );
  AOI22XL U4022 ( .A0(n3866), .A1(image_data[69]), .B0(n3867), .B1(
        image_data[197]), .Y(n4214) );
  NAND4XL U4023 ( .A(n4207), .B(n4206), .C(n4205), .D(n4204), .Y(n4208) );
  AOI22XL U4024 ( .A0(n3928), .A1(image_data[285]), .B0(n3929), .B1(
        image_data[413]), .Y(n4207) );
  AOI22XL U4025 ( .A0(n4702), .A1(image_data[349]), .B0(n3894), .B1(
        image_data[477]), .Y(n4206) );
  AOI22XL U4026 ( .A0(n3896), .A1(image_data[381]), .B0(n4670), .B1(
        image_data[509]), .Y(n4204) );
  NAND4XL U4027 ( .A(n4199), .B(n4198), .C(n4197), .D(n4196), .Y(n4210) );
  AOI22XL U4028 ( .A0(n3875), .A1(image_data[341]), .B0(n3876), .B1(
        image_data[469]), .Y(n4198) );
  AOI22XL U4029 ( .A0(n3877), .A1(image_data[309]), .B0(n3949), .B1(
        image_data[437]), .Y(n4197) );
  AOI22XL U4030 ( .A0(n3874), .A1(image_data[277]), .B0(n3948), .B1(
        image_data[405]), .Y(n4199) );
  NAND4XL U4031 ( .A(n4195), .B(n4194), .C(n4193), .D(n4192), .Y(n4211) );
  AOI22XL U4032 ( .A0(n3865), .A1(image_data[261]), .B0(n3941), .B1(
        image_data[389]), .Y(n4195) );
  AOI22XL U4033 ( .A0(n3866), .A1(image_data[325]), .B0(n3867), .B1(
        image_data[453]), .Y(n4194) );
  AOI22XL U4034 ( .A0(n3942), .A1(image_data[293]), .B0(n3943), .B1(
        image_data[421]), .Y(n4193) );
  AOI22XL U4035 ( .A0(n3884), .A1(image_data[341]), .B0(n3934), .B1(
        image_data[469]), .Y(n3987) );
  AOI22XL U4036 ( .A0(n3887), .A1(image_data[373]), .B0(n3936), .B1(
        image_data[501]), .Y(n3985) );
  AOI22XL U4037 ( .A0(n3888), .A1(image_data[309]), .B0(n4763), .B1(
        image_data[437]), .Y(n3986) );
  NAND4XL U4038 ( .A(n4016), .B(n4015), .C(n4014), .D(n4013), .Y(n4017) );
  AOI22XL U4039 ( .A0(n3876), .A1(image_data[29]), .B0(n3875), .B1(
        image_data[157]), .Y(n4016) );
  AOI22XL U4040 ( .A0(n3877), .A1(image_data[125]), .B0(n3949), .B1(
        image_data[253]), .Y(n4013) );
  AOI22XL U4041 ( .A0(n3874), .A1(image_data[93]), .B0(n3948), .B1(
        image_data[221]), .Y(n4015) );
  NAND4XL U4042 ( .A(n4012), .B(n4011), .C(n4010), .D(n4009), .Y(n4018) );
  AOI22XL U4043 ( .A0(n3867), .A1(image_data[13]), .B0(n3866), .B1(
        image_data[141]), .Y(n4012) );
  AOI22XL U4044 ( .A0(n3865), .A1(image_data[77]), .B0(n3941), .B1(
        image_data[205]), .Y(n4011) );
  AOI22XL U4045 ( .A0(n3942), .A1(image_data[109]), .B0(n3943), .B1(
        image_data[237]), .Y(n4009) );
  NAND4XL U4046 ( .A(n4004), .B(n4003), .C(n4002), .D(n4001), .Y(n4020) );
  AOI22XL U4047 ( .A0(n3364), .A1(image_data[5]), .B0(n4681), .B1(
        image_data[133]), .Y(n4004) );
  AOI22XL U4048 ( .A0(n3897), .A1(image_data[69]), .B0(n3896), .B1(
        image_data[197]), .Y(n4003) );
  AOI22XL U4049 ( .A0(n3928), .A1(image_data[101]), .B0(n3929), .B1(
        image_data[229]), .Y(n4001) );
  NAND4XL U4050 ( .A(n4008), .B(n4007), .C(n4006), .D(n4005), .Y(n4019) );
  AOI22XL U4051 ( .A0(n3886), .A1(image_data[21]), .B0(n3885), .B1(
        image_data[149]), .Y(n4008) );
  AOI22XL U4052 ( .A0(n3888), .A1(image_data[53]), .B0(n4763), .B1(
        image_data[181]), .Y(n4006) );
  AOI22XL U4053 ( .A0(n3887), .A1(image_data[117]), .B0(n3936), .B1(
        image_data[245]), .Y(n4005) );
  NAND4XL U4054 ( .A(n3996), .B(n3995), .C(n3994), .D(n3993), .Y(n3997) );
  AOI22XL U4055 ( .A0(n3876), .A1(image_data[285]), .B0(n3875), .B1(
        image_data[413]), .Y(n3996) );
  AOI22XL U4056 ( .A0(n3877), .A1(image_data[381]), .B0(n3949), .B1(
        image_data[509]), .Y(n3993) );
  AOI22XL U4057 ( .A0(n3874), .A1(image_data[349]), .B0(n3948), .B1(
        image_data[477]), .Y(n3995) );
  NAND4XL U4058 ( .A(n3992), .B(n3991), .C(n3990), .D(n3989), .Y(n3998) );
  AOI22XL U4059 ( .A0(n3867), .A1(image_data[269]), .B0(n3866), .B1(
        image_data[397]), .Y(n3992) );
  AOI22XL U4060 ( .A0(n3865), .A1(image_data[333]), .B0(n3941), .B1(
        image_data[461]), .Y(n3991) );
  AOI22XL U4061 ( .A0(n3942), .A1(image_data[365]), .B0(n3943), .B1(
        image_data[493]), .Y(n3989) );
  NAND4XL U4062 ( .A(n3984), .B(n3983), .C(n3982), .D(n3981), .Y(n4000) );
  AOI22XL U4063 ( .A0(n3928), .A1(image_data[357]), .B0(n3929), .B1(
        image_data[485]), .Y(n3981) );
  AOI22XL U4064 ( .A0(n3897), .A1(image_data[325]), .B0(n3896), .B1(
        image_data[453]), .Y(n3983) );
  AOI22XL U4065 ( .A0(n3894), .A1(image_data[293]), .B0(n3893), .B1(
        image_data[421]), .Y(n3982) );
  AOI22XL U4066 ( .A0(n3942), .A1(image_data[294]), .B0(n3943), .B1(
        image_data[422]), .Y(n4319) );
  AOI22XL U4067 ( .A0(n3865), .A1(image_data[262]), .B0(n3941), .B1(
        image_data[390]), .Y(n4321) );
  AOI22XL U4068 ( .A0(n4714), .A1(image_data[358]), .B0(n3869), .B1(
        image_data[486]), .Y(n4318) );
  AOI22XL U4069 ( .A0(n3866), .A1(image_data[326]), .B0(n3867), .B1(
        image_data[454]), .Y(n4320) );
  NAND4XL U4070 ( .A(n4353), .B(n4352), .C(n4351), .D(n4350), .Y(n4354) );
  AOI22XL U4071 ( .A0(n3896), .A1(image_data[126]), .B0(n3897), .B1(
        image_data[254]), .Y(n4350) );
  AOI22XL U4072 ( .A0(n3928), .A1(image_data[30]), .B0(n3929), .B1(
        image_data[158]), .Y(n4353) );
  AOI22XL U4073 ( .A0(n3893), .A1(image_data[94]), .B0(n3894), .B1(
        image_data[222]), .Y(n4352) );
  NAND4XL U4074 ( .A(n4349), .B(n4348), .C(n4347), .D(n4346), .Y(n4355) );
  AOI22XL U4075 ( .A0(n3885), .A1(image_data[78]), .B0(n3886), .B1(
        image_data[206]), .Y(n4348) );
  AOI22XL U4076 ( .A0(n4763), .A1(image_data[110]), .B0(n3888), .B1(
        image_data[238]), .Y(n4346) );
  AOI22XL U4077 ( .A0(n3887), .A1(image_data[46]), .B0(n3936), .B1(
        image_data[174]), .Y(n4347) );
  NAND4XL U4078 ( .A(n4345), .B(n4344), .C(n4343), .D(n4342), .Y(n4356) );
  AOI22XL U4079 ( .A0(n4719), .A1(image_data[86]), .B0(n3876), .B1(
        image_data[214]), .Y(n4344) );
  AOI22XL U4080 ( .A0(n4721), .A1(image_data[118]), .B0(n3879), .B1(
        image_data[246]), .Y(n4342) );
  AOI22XL U4081 ( .A0(n3877), .A1(image_data[54]), .B0(n3949), .B1(
        image_data[182]), .Y(n4343) );
  NAND4XL U4082 ( .A(n4341), .B(n4340), .C(n4339), .D(n4338), .Y(n4357) );
  AOI22XL U4083 ( .A0(n4714), .A1(image_data[102]), .B0(n3869), .B1(
        image_data[230]), .Y(n4338) );
  AOI22XL U4084 ( .A0(n3866), .A1(image_data[70]), .B0(n3867), .B1(
        image_data[198]), .Y(n4340) );
  AOI22XL U4085 ( .A0(n3865), .A1(image_data[6]), .B0(n3941), .B1(
        image_data[134]), .Y(n4341) );
  NAND4XL U4086 ( .A(n4333), .B(n4332), .C(n4331), .D(n4330), .Y(n4334) );
  AOI22XL U4087 ( .A0(n3896), .A1(image_data[382]), .B0(n3897), .B1(
        image_data[510]), .Y(n4330) );
  AOI22XL U4088 ( .A0(n4702), .A1(image_data[350]), .B0(n3894), .B1(
        image_data[478]), .Y(n4332) );
  AOI22XL U4089 ( .A0(n3928), .A1(image_data[286]), .B0(n3929), .B1(
        image_data[414]), .Y(n4333) );
  NAND4XL U4090 ( .A(n4329), .B(n4328), .C(n4327), .D(n4326), .Y(n4335) );
  AOI22XL U4091 ( .A0(n4707), .A1(image_data[334]), .B0(n3886), .B1(
        image_data[462]), .Y(n4328) );
  AOI22XL U4092 ( .A0(n4763), .A1(image_data[366]), .B0(n3888), .B1(
        image_data[494]), .Y(n4326) );
  AOI22XL U4093 ( .A0(n3887), .A1(image_data[302]), .B0(n3936), .B1(
        image_data[430]), .Y(n4327) );
  NAND4XL U4094 ( .A(n4325), .B(n4324), .C(n4323), .D(n4322), .Y(n4336) );
  AOI22XL U4095 ( .A0(n4719), .A1(image_data[342]), .B0(n3876), .B1(
        image_data[470]), .Y(n4324) );
  AOI22XL U4096 ( .A0(n4721), .A1(image_data[374]), .B0(n3879), .B1(
        image_data[502]), .Y(n4322) );
  AOI22XL U4097 ( .A0(n3877), .A1(image_data[310]), .B0(n3949), .B1(
        image_data[438]), .Y(n4323) );
  AOI22XL U4098 ( .A0(n3942), .A1(image_data[290]), .B0(n3943), .B1(
        image_data[418]), .Y(n3871) );
  AOI22XL U4099 ( .A0(n3865), .A1(image_data[258]), .B0(n3941), .B1(
        image_data[386]), .Y(n3873) );
  AOI22XL U4100 ( .A0(n4714), .A1(image_data[354]), .B0(n3869), .B1(
        image_data[482]), .Y(n3870) );
  AOI22XL U4101 ( .A0(n3866), .A1(image_data[322]), .B0(n3867), .B1(
        image_data[450]), .Y(n3872) );
  NAND4XL U4102 ( .A(n3921), .B(n3920), .C(n3919), .D(n3918), .Y(n3922) );
  AOI22XL U4103 ( .A0(n3896), .A1(image_data[122]), .B0(n3897), .B1(
        image_data[250]), .Y(n3918) );
  AOI22XL U4104 ( .A0(n3928), .A1(image_data[26]), .B0(n3929), .B1(
        image_data[154]), .Y(n3921) );
  AOI22XL U4105 ( .A0(n3893), .A1(image_data[90]), .B0(n3894), .B1(
        image_data[218]), .Y(n3920) );
  NAND4XL U4106 ( .A(n3917), .B(n3916), .C(n3915), .D(n3914), .Y(n3923) );
  AOI22XL U4107 ( .A0(n3885), .A1(image_data[74]), .B0(n3886), .B1(
        image_data[202]), .Y(n3916) );
  AOI22XL U4108 ( .A0(n3935), .A1(image_data[106]), .B0(n3888), .B1(
        image_data[234]), .Y(n3914) );
  AOI22XL U4109 ( .A0(n3884), .A1(image_data[10]), .B0(n3934), .B1(
        image_data[138]), .Y(n3917) );
  NAND4XL U4110 ( .A(n3913), .B(n3912), .C(n3911), .D(n3910), .Y(n3924) );
  AOI22XL U4111 ( .A0(n3875), .A1(image_data[82]), .B0(n3876), .B1(
        image_data[210]), .Y(n3912) );
  AOI22XL U4112 ( .A0(n3877), .A1(image_data[50]), .B0(n3949), .B1(
        image_data[178]), .Y(n3911) );
  AOI22XL U4113 ( .A0(n3874), .A1(image_data[18]), .B0(n3948), .B1(
        image_data[146]), .Y(n3913) );
  NAND4XL U4114 ( .A(n3909), .B(n3908), .C(n3907), .D(n3906), .Y(n3925) );
  AOI22XL U4115 ( .A0(n3866), .A1(image_data[66]), .B0(n3867), .B1(
        image_data[194]), .Y(n3908) );
  AOI22XL U4116 ( .A0(n4714), .A1(image_data[98]), .B0(n3869), .B1(
        image_data[226]), .Y(n3906) );
  AOI22XL U4117 ( .A0(n3865), .A1(image_data[2]), .B0(n3941), .B1(
        image_data[130]), .Y(n3909) );
  NAND4XL U4118 ( .A(n3901), .B(n3900), .C(n3899), .D(n3898), .Y(n3902) );
  AOI22XL U4119 ( .A0(n4702), .A1(image_data[346]), .B0(n3894), .B1(
        image_data[474]), .Y(n3900) );
  AOI22XL U4120 ( .A0(n3896), .A1(image_data[378]), .B0(n3897), .B1(
        image_data[506]), .Y(n3898) );
  AOI22XL U4121 ( .A0(n3928), .A1(image_data[282]), .B0(n3929), .B1(
        image_data[410]), .Y(n3901) );
  NAND4XL U4122 ( .A(n3892), .B(n3891), .C(n3890), .D(n3889), .Y(n3903) );
  AOI22XL U4123 ( .A0(n3885), .A1(image_data[330]), .B0(n3886), .B1(
        image_data[458]), .Y(n3891) );
  AOI22XL U4124 ( .A0(n3935), .A1(image_data[362]), .B0(n3888), .B1(
        image_data[490]), .Y(n3889) );
  AOI22XL U4125 ( .A0(n3884), .A1(image_data[266]), .B0(n3934), .B1(
        image_data[394]), .Y(n3892) );
  NAND4XL U4126 ( .A(n3883), .B(n3882), .C(n3881), .D(n3880), .Y(n3904) );
  AOI22XL U4127 ( .A0(n3875), .A1(image_data[338]), .B0(n3876), .B1(
        image_data[466]), .Y(n3882) );
  AOI22XL U4128 ( .A0(n4721), .A1(image_data[370]), .B0(n3879), .B1(
        image_data[498]), .Y(n3880) );
  AOI22XL U4129 ( .A0(n3877), .A1(image_data[306]), .B0(n3949), .B1(
        image_data[434]), .Y(n3881) );
  AOI22XL U4130 ( .A0(n4714), .A1(image_data[359]), .B0(n3869), .B1(
        image_data[487]), .Y(n4360) );
  AOI22XL U4131 ( .A0(n3942), .A1(image_data[295]), .B0(n3943), .B1(
        image_data[423]), .Y(n4361) );
  NAND4XL U4132 ( .A(n4395), .B(n4394), .C(n4393), .D(n4392), .Y(n4396) );
  AOI22XL U4133 ( .A0(n4681), .A1(image_data[63]), .B0(n3364), .B1(
        image_data[191]), .Y(n4393) );
  AOI22XL U4134 ( .A0(n3928), .A1(image_data[31]), .B0(n3929), .B1(
        image_data[159]), .Y(n4395) );
  AOI22XL U4135 ( .A0(n4702), .A1(image_data[95]), .B0(n3894), .B1(
        image_data[223]), .Y(n4394) );
  NAND4XL U4136 ( .A(n4391), .B(n4390), .C(n4389), .D(n4388), .Y(n4397) );
  AOI22XL U4137 ( .A0(n4707), .A1(image_data[79]), .B0(n3886), .B1(
        image_data[207]), .Y(n4390) );
  AOI22XL U4138 ( .A0(n3887), .A1(image_data[47]), .B0(n3936), .B1(
        image_data[175]), .Y(n4389) );
  AOI22XL U4139 ( .A0(n3884), .A1(image_data[15]), .B0(n3934), .B1(
        image_data[143]), .Y(n4391) );
  NAND4XL U4140 ( .A(n4387), .B(n4386), .C(n4385), .D(n4384), .Y(n4398) );
  AOI22XL U4141 ( .A0(n4719), .A1(image_data[87]), .B0(n3876), .B1(
        image_data[215]), .Y(n4386) );
  AOI22XL U4142 ( .A0(n3877), .A1(image_data[55]), .B0(n3949), .B1(
        image_data[183]), .Y(n4385) );
  AOI22XL U4143 ( .A0(n3874), .A1(image_data[23]), .B0(n3948), .B1(
        image_data[151]), .Y(n4387) );
  NAND4XL U4144 ( .A(n4383), .B(n4382), .C(n4381), .D(n4380), .Y(n4399) );
  AOI22XL U4145 ( .A0(n3865), .A1(image_data[7]), .B0(n3941), .B1(
        image_data[135]), .Y(n4383) );
  AOI22XL U4146 ( .A0(n3866), .A1(image_data[71]), .B0(n3867), .B1(
        image_data[199]), .Y(n4382) );
  AOI22XL U4147 ( .A0(n3942), .A1(image_data[39]), .B0(n3943), .B1(
        image_data[167]), .Y(n4381) );
  NAND4XL U4148 ( .A(n4375), .B(n4374), .C(n4373), .D(n4372), .Y(n4376) );
  AOI22XL U4149 ( .A0(n4681), .A1(image_data[319]), .B0(n3364), .B1(
        image_data[447]), .Y(n4373) );
  AOI22XL U4150 ( .A0(n3928), .A1(image_data[287]), .B0(n3929), .B1(
        image_data[415]), .Y(n4375) );
  AOI22XL U4151 ( .A0(n3896), .A1(image_data[383]), .B0(n3897), .B1(
        image_data[511]), .Y(n4372) );
  NAND4XL U4152 ( .A(n4371), .B(n4370), .C(n4369), .D(n4368), .Y(n4377) );
  AOI22XL U4153 ( .A0(n4707), .A1(image_data[335]), .B0(n3886), .B1(
        image_data[463]), .Y(n4370) );
  AOI22XL U4154 ( .A0(n3887), .A1(image_data[303]), .B0(n3936), .B1(
        image_data[431]), .Y(n4369) );
  AOI22XL U4155 ( .A0(n3884), .A1(image_data[271]), .B0(n3934), .B1(
        image_data[399]), .Y(n4371) );
  NAND4XL U4156 ( .A(n4367), .B(n4366), .C(n4365), .D(n4364), .Y(n4378) );
  AOI22XL U4157 ( .A0(n4719), .A1(image_data[343]), .B0(n3876), .B1(
        image_data[471]), .Y(n4366) );
  AOI22XL U4158 ( .A0(n3877), .A1(image_data[311]), .B0(n3949), .B1(
        image_data[439]), .Y(n4365) );
  AOI22XL U4159 ( .A0(n3874), .A1(image_data[279]), .B0(n3948), .B1(
        image_data[407]), .Y(n4367) );
  INVX1 U4160 ( .A(n6820), .Y(n6802) );
  NOR4XL U4161 ( .A(n4938), .B(n4937), .C(n4936), .D(n4935), .Y(n4961) );
  NOR4XL U4162 ( .A(n4958), .B(n4957), .C(n4956), .D(n4955), .Y(n4960) );
  NAND4XL U4163 ( .A(n4926), .B(n4925), .C(n4924), .D(n4923), .Y(n4937) );
  NOR4XL U4164 ( .A(n4657), .B(n4656), .C(n4655), .D(n4654), .Y(n4680) );
  NOR4XL U4165 ( .A(n4678), .B(n4677), .C(n4676), .D(n4675), .Y(n4679) );
  NAND4XL U4166 ( .A(n4649), .B(n4648), .C(n4647), .D(n4646), .Y(n4655) );
  NOR4XL U4167 ( .A(n4896), .B(n4895), .C(n4894), .D(n4893), .Y(n4918) );
  NOR4XL U4168 ( .A(n4916), .B(n4915), .C(n4914), .D(n4913), .Y(n4917) );
  NAND4XL U4169 ( .A(n4892), .B(n4891), .C(n4890), .D(n4889), .Y(n4893) );
  NOR4XL U4170 ( .A(n4752), .B(n4751), .C(n4750), .D(n4749), .Y(n4779) );
  NOR4XL U4171 ( .A(n4776), .B(n4775), .C(n4774), .D(n4773), .Y(n4778) );
  NAND4XL U4172 ( .A(n4744), .B(n4743), .C(n4742), .D(n4741), .Y(n4750) );
  NOR4XL U4173 ( .A(n4847), .B(n4846), .C(n4845), .D(n4844), .Y(n4870) );
  NOR4XL U4174 ( .A(n4867), .B(n4866), .C(n4865), .D(n4864), .Y(n4869) );
  NOR4XL U4175 ( .A(n4701), .B(n4700), .C(n4699), .D(n4698), .Y(n4732) );
  NOR4XL U4176 ( .A(n4730), .B(n4729), .C(n4728), .D(n4727), .Y(n4731) );
  NAND4XL U4177 ( .A(n4689), .B(n4688), .C(n4687), .D(n4686), .Y(n4700) );
  AOI22XL U4178 ( .A0(n6498), .A1(n5854), .B0(n5853), .B1(n6495), .Y(n5900) );
  AOI22XL U4179 ( .A0(n6574), .A1(n5896), .B0(n5895), .B1(n6571), .Y(n5899) );
  NOR4XL U4180 ( .A(n5832), .B(n5831), .C(n5830), .D(n5829), .Y(n5854) );
  AOI22XL U4181 ( .A0(n6498), .A1(n5751), .B0(n5750), .B1(n6495), .Y(n5797) );
  AOI22XL U4182 ( .A0(n6574), .A1(n5793), .B0(n5792), .B1(n6571), .Y(n5796) );
  NOR4XL U4183 ( .A(n5729), .B(n5728), .C(n5727), .D(n5726), .Y(n5751) );
  NOR4XL U4184 ( .A(n4512), .B(n4511), .C(n4510), .D(n4509), .Y(n4534) );
  NOR4XL U4185 ( .A(n4532), .B(n4531), .C(n4530), .D(n4529), .Y(n4533) );
  NAND4XL U4186 ( .A(n4500), .B(n4499), .C(n4498), .D(n4497), .Y(n4511) );
  AOI22X2 U4187 ( .A0(n5165), .A1(n3559), .B0(n3558), .B1(n4777), .Y(N2781) );
  NAND4XL U4188 ( .A(n3521), .B(n3520), .C(n3519), .D(n3518), .Y(n3537) );
  NAND4XL U4189 ( .A(n4245), .B(n4244), .C(n4243), .D(n4242), .Y(n4251) );
  NAND4XL U4190 ( .A(n4157), .B(n4156), .C(n4155), .D(n4154), .Y(n4168) );
  NOR4XL U4191 ( .A(n4127), .B(n4126), .C(n4125), .D(n4124), .Y(n4149) );
  NOR4XL U4192 ( .A(n4147), .B(n4146), .C(n4145), .D(n4144), .Y(n4148) );
  NAND4XL U4193 ( .A(n4115), .B(n4114), .C(n4113), .D(n4112), .Y(n4126) );
  INVXL U4194 ( .A(N2759), .Y(n6173) );
  AOI22X2 U4195 ( .A0(n3450), .A1(n3601), .B0(n3600), .B1(n4959), .Y(N2755) );
  NAND4XL U4196 ( .A(n3567), .B(n3566), .C(n3565), .D(n3564), .Y(n3578) );
  AOI22X2 U4197 ( .A0(n5165), .A1(n3643), .B0(n3642), .B1(n4777), .Y(N2779) );
  NOR4X1 U4198 ( .A(n3621), .B(n3620), .C(n3619), .D(n3618), .Y(n3643) );
  NOR4X1 U4199 ( .A(n3641), .B(n3640), .C(n3639), .D(n3638), .Y(n3642) );
  NAND4XL U4200 ( .A(n3605), .B(n3604), .C(n3603), .D(n3602), .Y(n3621) );
  NAND4XL U4201 ( .A(n5518), .B(n5517), .C(n5516), .D(n5515), .Y(n5519) );
  AOI22XL U4202 ( .A0(n5584), .A1(image_data[88]), .B0(n5583), .B1(
        image_data[216]), .Y(n5517) );
  AOI22XL U4203 ( .A0(n5586), .A1(image_data[56]), .B0(n5585), .B1(
        image_data[184]), .Y(n5516) );
  AOI22XL U4204 ( .A0(n5588), .A1(image_data[120]), .B0(n5587), .B1(
        image_data[248]), .Y(n5515) );
  NAND4XL U4205 ( .A(n5514), .B(n5513), .C(n5512), .D(n5511), .Y(n5520) );
  AOI22XL U4206 ( .A0(n5572), .A1(image_data[72]), .B0(n5571), .B1(
        image_data[200]), .Y(n5513) );
  AOI22XL U4207 ( .A0(n5574), .A1(image_data[40]), .B0(n5573), .B1(
        image_data[168]), .Y(n5512) );
  AOI22XL U4208 ( .A0(n5576), .A1(image_data[104]), .B0(n5575), .B1(
        image_data[232]), .Y(n5511) );
  NAND4XL U4209 ( .A(n5510), .B(n5509), .C(n5508), .D(n5507), .Y(n5521) );
  AOI22XL U4210 ( .A0(n5560), .A1(image_data[80]), .B0(n5559), .B1(
        image_data[208]), .Y(n5509) );
  AOI22XL U4211 ( .A0(n5562), .A1(image_data[48]), .B0(n5561), .B1(
        image_data[176]), .Y(n5508) );
  AOI22XL U4212 ( .A0(n5564), .A1(image_data[112]), .B0(n5563), .B1(
        image_data[240]), .Y(n5507) );
  NAND4XL U4213 ( .A(n5498), .B(n5497), .C(n5496), .D(n5495), .Y(n5499) );
  AOI22XL U4214 ( .A0(n5584), .A1(image_data[344]), .B0(n5583), .B1(
        image_data[472]), .Y(n5497) );
  AOI22XL U4215 ( .A0(n5586), .A1(image_data[312]), .B0(n5585), .B1(
        image_data[440]), .Y(n5496) );
  AOI22XL U4216 ( .A0(n5588), .A1(image_data[376]), .B0(n5587), .B1(
        image_data[504]), .Y(n5495) );
  NAND4XL U4217 ( .A(n5494), .B(n5493), .C(n5492), .D(n5491), .Y(n5500) );
  AOI22XL U4218 ( .A0(n5572), .A1(image_data[328]), .B0(n5571), .B1(
        image_data[456]), .Y(n5493) );
  AOI22XL U4219 ( .A0(n5574), .A1(image_data[296]), .B0(n5573), .B1(
        image_data[424]), .Y(n5492) );
  AOI22XL U4220 ( .A0(n5576), .A1(image_data[360]), .B0(n5575), .B1(
        image_data[488]), .Y(n5491) );
  NAND4XL U4221 ( .A(n5434), .B(n5433), .C(n5432), .D(n5431), .Y(n5435) );
  AOI22XL U4222 ( .A0(n5584), .A1(image_data[89]), .B0(n5583), .B1(
        image_data[217]), .Y(n5433) );
  AOI22XL U4223 ( .A0(n5586), .A1(image_data[57]), .B0(n5585), .B1(
        image_data[185]), .Y(n5432) );
  AOI22XL U4224 ( .A0(n5588), .A1(image_data[121]), .B0(n5587), .B1(
        image_data[249]), .Y(n5431) );
  NAND4XL U4225 ( .A(n5430), .B(n5429), .C(n5428), .D(n5427), .Y(n5436) );
  AOI22XL U4226 ( .A0(n5572), .A1(image_data[73]), .B0(n5571), .B1(
        image_data[201]), .Y(n5429) );
  AOI22XL U4227 ( .A0(n5574), .A1(image_data[41]), .B0(n5573), .B1(
        image_data[169]), .Y(n5428) );
  AOI22XL U4228 ( .A0(n5576), .A1(image_data[105]), .B0(n5575), .B1(
        image_data[233]), .Y(n5427) );
  NAND4XL U4229 ( .A(n5426), .B(n5425), .C(n5424), .D(n5423), .Y(n5437) );
  AOI22XL U4230 ( .A0(n5560), .A1(image_data[81]), .B0(n5559), .B1(
        image_data[209]), .Y(n5425) );
  AOI22XL U4231 ( .A0(n5562), .A1(image_data[49]), .B0(n5561), .B1(
        image_data[177]), .Y(n5424) );
  AOI22XL U4232 ( .A0(n5564), .A1(image_data[113]), .B0(n5563), .B1(
        image_data[241]), .Y(n5423) );
  NAND4XL U4233 ( .A(n5414), .B(n5413), .C(n5412), .D(n5411), .Y(n5415) );
  AOI22XL U4234 ( .A0(n5584), .A1(image_data[345]), .B0(n5583), .B1(
        image_data[473]), .Y(n5413) );
  AOI22XL U4235 ( .A0(n5586), .A1(image_data[313]), .B0(n5585), .B1(
        image_data[441]), .Y(n5412) );
  AOI22XL U4236 ( .A0(n5588), .A1(image_data[377]), .B0(n5587), .B1(
        image_data[505]), .Y(n5411) );
  NAND4XL U4237 ( .A(n5410), .B(n5409), .C(n5408), .D(n5407), .Y(n5416) );
  AOI22XL U4238 ( .A0(n5572), .A1(image_data[329]), .B0(n5571), .B1(
        image_data[457]), .Y(n5409) );
  AOI22XL U4239 ( .A0(n5574), .A1(image_data[297]), .B0(n5573), .B1(
        image_data[425]), .Y(n5408) );
  AOI22XL U4240 ( .A0(n5576), .A1(image_data[361]), .B0(n5575), .B1(
        image_data[489]), .Y(n5407) );
  NAND4XL U4241 ( .A(n4580), .B(n4579), .C(n4578), .D(n4577), .Y(n4581) );
  AOI22XL U4242 ( .A0(n5584), .A1(image_data[90]), .B0(n5583), .B1(
        image_data[218]), .Y(n4579) );
  AOI22XL U4243 ( .A0(n5586), .A1(image_data[58]), .B0(n5585), .B1(
        image_data[186]), .Y(n4578) );
  AOI22XL U4244 ( .A0(n5588), .A1(image_data[122]), .B0(n5587), .B1(
        image_data[250]), .Y(n4577) );
  NAND4XL U4245 ( .A(n4576), .B(n4575), .C(n4574), .D(n4573), .Y(n4582) );
  AOI22XL U4246 ( .A0(n5572), .A1(image_data[74]), .B0(n5571), .B1(
        image_data[202]), .Y(n4575) );
  AOI22XL U4247 ( .A0(n5574), .A1(image_data[42]), .B0(n5573), .B1(
        image_data[170]), .Y(n4574) );
  AOI22XL U4248 ( .A0(n5576), .A1(image_data[106]), .B0(n5575), .B1(
        image_data[234]), .Y(n4573) );
  NAND4XL U4249 ( .A(n4572), .B(n4571), .C(n4570), .D(n4569), .Y(n4583) );
  AOI22XL U4250 ( .A0(n5560), .A1(image_data[82]), .B0(n5559), .B1(
        image_data[210]), .Y(n4571) );
  AOI22XL U4251 ( .A0(n5562), .A1(image_data[50]), .B0(n5561), .B1(
        image_data[178]), .Y(n4570) );
  AOI22XL U4252 ( .A0(n5564), .A1(image_data[114]), .B0(n5563), .B1(
        image_data[242]), .Y(n4569) );
  NAND4XL U4253 ( .A(n4560), .B(n4559), .C(n4558), .D(n4557), .Y(n4561) );
  AOI22XL U4254 ( .A0(n5584), .A1(image_data[346]), .B0(n5583), .B1(
        image_data[474]), .Y(n4559) );
  AOI22XL U4255 ( .A0(n5586), .A1(image_data[314]), .B0(n5585), .B1(
        image_data[442]), .Y(n4558) );
  AOI22XL U4256 ( .A0(n5588), .A1(image_data[378]), .B0(n5587), .B1(
        image_data[506]), .Y(n4557) );
  NAND4XL U4257 ( .A(n4548), .B(n4547), .C(n4546), .D(n4545), .Y(n4562) );
  AOI22XL U4258 ( .A0(n5572), .A1(image_data[330]), .B0(n5571), .B1(
        image_data[458]), .Y(n4547) );
  AOI22XL U4259 ( .A0(n5574), .A1(image_data[298]), .B0(n5573), .B1(
        image_data[426]), .Y(n4546) );
  AOI22XL U4260 ( .A0(n5576), .A1(image_data[362]), .B0(n5575), .B1(
        image_data[490]), .Y(n4545) );
  NAND4XL U4261 ( .A(n5592), .B(n5591), .C(n5590), .D(n5589), .Y(n5593) );
  AOI22XL U4262 ( .A0(n5584), .A1(image_data[91]), .B0(n5583), .B1(
        image_data[219]), .Y(n5591) );
  AOI22XL U4263 ( .A0(n5586), .A1(image_data[59]), .B0(n5585), .B1(
        image_data[187]), .Y(n5590) );
  AOI22XL U4264 ( .A0(n5588), .A1(image_data[123]), .B0(n5587), .B1(
        image_data[251]), .Y(n5589) );
  NAND4XL U4265 ( .A(n5580), .B(n5579), .C(n5578), .D(n5577), .Y(n5594) );
  AOI22XL U4266 ( .A0(n5572), .A1(image_data[75]), .B0(n5571), .B1(
        image_data[203]), .Y(n5579) );
  AOI22XL U4267 ( .A0(n5574), .A1(image_data[43]), .B0(n5573), .B1(
        image_data[171]), .Y(n5578) );
  AOI22XL U4268 ( .A0(n5576), .A1(image_data[107]), .B0(n5575), .B1(
        image_data[235]), .Y(n5577) );
  NAND4XL U4269 ( .A(n5568), .B(n5567), .C(n5566), .D(n5565), .Y(n5595) );
  AOI22XL U4270 ( .A0(n5560), .A1(image_data[83]), .B0(n5559), .B1(
        image_data[211]), .Y(n5567) );
  AOI22XL U4271 ( .A0(n5562), .A1(image_data[51]), .B0(n5561), .B1(
        image_data[179]), .Y(n5566) );
  AOI22XL U4272 ( .A0(n5564), .A1(image_data[115]), .B0(n5563), .B1(
        image_data[243]), .Y(n5565) );
  NAND4XL U4273 ( .A(n5540), .B(n5539), .C(n5538), .D(n5537), .Y(n5541) );
  AOI22XL U4274 ( .A0(n5584), .A1(image_data[347]), .B0(n5583), .B1(
        image_data[475]), .Y(n5539) );
  AOI22XL U4275 ( .A0(n5586), .A1(image_data[315]), .B0(n5585), .B1(
        image_data[443]), .Y(n5538) );
  AOI22XL U4276 ( .A0(n5588), .A1(image_data[379]), .B0(n5587), .B1(
        image_data[507]), .Y(n5537) );
  NAND4XL U4277 ( .A(n5536), .B(n5535), .C(n5534), .D(n5533), .Y(n5542) );
  AOI22XL U4278 ( .A0(n5572), .A1(image_data[331]), .B0(n5571), .B1(
        image_data[459]), .Y(n5535) );
  AOI22XL U4279 ( .A0(n5574), .A1(image_data[299]), .B0(n5573), .B1(
        image_data[427]), .Y(n5534) );
  AOI22XL U4280 ( .A0(n5576), .A1(image_data[363]), .B0(n5575), .B1(
        image_data[491]), .Y(n5533) );
  NAND4XL U4281 ( .A(n5476), .B(n5475), .C(n5474), .D(n5473), .Y(n5477) );
  AOI22XL U4282 ( .A0(n5584), .A1(image_data[92]), .B0(n5583), .B1(
        image_data[220]), .Y(n5475) );
  AOI22XL U4283 ( .A0(n5586), .A1(image_data[60]), .B0(n5585), .B1(
        image_data[188]), .Y(n5474) );
  AOI22XL U4284 ( .A0(n5588), .A1(image_data[124]), .B0(n5587), .B1(
        image_data[252]), .Y(n5473) );
  NAND4XL U4285 ( .A(n5472), .B(n5471), .C(n5470), .D(n5469), .Y(n5478) );
  AOI22XL U4286 ( .A0(n5572), .A1(image_data[76]), .B0(n5571), .B1(
        image_data[204]), .Y(n5471) );
  AOI22XL U4287 ( .A0(n5574), .A1(image_data[44]), .B0(n5573), .B1(
        image_data[172]), .Y(n5470) );
  AOI22XL U4288 ( .A0(n5576), .A1(image_data[108]), .B0(n5575), .B1(
        image_data[236]), .Y(n5469) );
  NAND4XL U4289 ( .A(n5468), .B(n5467), .C(n5466), .D(n5465), .Y(n5479) );
  AOI22XL U4290 ( .A0(n5560), .A1(image_data[84]), .B0(n5559), .B1(
        image_data[212]), .Y(n5467) );
  AOI22XL U4291 ( .A0(n5562), .A1(image_data[52]), .B0(n5561), .B1(
        image_data[180]), .Y(n5466) );
  AOI22XL U4292 ( .A0(n5564), .A1(image_data[116]), .B0(n5563), .B1(
        image_data[244]), .Y(n5465) );
  NAND4XL U4293 ( .A(n5456), .B(n5455), .C(n5454), .D(n5453), .Y(n5457) );
  AOI22XL U4294 ( .A0(n5584), .A1(image_data[348]), .B0(n5583), .B1(
        image_data[476]), .Y(n5455) );
  AOI22XL U4295 ( .A0(n5586), .A1(image_data[316]), .B0(n5585), .B1(
        image_data[444]), .Y(n5454) );
  AOI22XL U4296 ( .A0(n5588), .A1(image_data[380]), .B0(n5587), .B1(
        image_data[508]), .Y(n5453) );
  NAND4XL U4297 ( .A(n5452), .B(n5451), .C(n5450), .D(n5449), .Y(n5458) );
  AOI22XL U4298 ( .A0(n5572), .A1(image_data[332]), .B0(n5571), .B1(
        image_data[460]), .Y(n5451) );
  AOI22XL U4299 ( .A0(n5574), .A1(image_data[300]), .B0(n5573), .B1(
        image_data[428]), .Y(n5450) );
  AOI22XL U4300 ( .A0(n5576), .A1(image_data[364]), .B0(n5575), .B1(
        image_data[492]), .Y(n5449) );
  NAND4XL U4301 ( .A(n5392), .B(n5391), .C(n5390), .D(n5389), .Y(n5393) );
  AOI22XL U4302 ( .A0(n5584), .A1(image_data[93]), .B0(n5583), .B1(
        image_data[221]), .Y(n5391) );
  AOI22XL U4303 ( .A0(n5586), .A1(image_data[61]), .B0(n5585), .B1(
        image_data[189]), .Y(n5390) );
  AOI22XL U4304 ( .A0(n5588), .A1(image_data[125]), .B0(n5587), .B1(
        image_data[253]), .Y(n5389) );
  NAND4XL U4305 ( .A(n5388), .B(n5387), .C(n5386), .D(n5385), .Y(n5394) );
  AOI22XL U4306 ( .A0(n5572), .A1(image_data[77]), .B0(n5571), .B1(
        image_data[205]), .Y(n5387) );
  AOI22XL U4307 ( .A0(n5574), .A1(image_data[45]), .B0(n5573), .B1(
        image_data[173]), .Y(n5386) );
  AOI22XL U4308 ( .A0(n5576), .A1(image_data[109]), .B0(n5575), .B1(
        image_data[237]), .Y(n5385) );
  NAND4XL U4309 ( .A(n5384), .B(n5383), .C(n5382), .D(n5381), .Y(n5395) );
  AOI22XL U4310 ( .A0(n5560), .A1(image_data[85]), .B0(n5559), .B1(
        image_data[213]), .Y(n5383) );
  AOI22XL U4311 ( .A0(n5562), .A1(image_data[53]), .B0(n5561), .B1(
        image_data[181]), .Y(n5382) );
  AOI22XL U4312 ( .A0(n5564), .A1(image_data[117]), .B0(n5563), .B1(
        image_data[245]), .Y(n5381) );
  NAND4XL U4313 ( .A(n5372), .B(n5371), .C(n5370), .D(n5369), .Y(n5373) );
  AOI22XL U4314 ( .A0(n5584), .A1(image_data[349]), .B0(n5583), .B1(
        image_data[477]), .Y(n5371) );
  AOI22XL U4315 ( .A0(n5586), .A1(image_data[317]), .B0(n5585), .B1(
        image_data[445]), .Y(n5370) );
  AOI22XL U4316 ( .A0(n5588), .A1(image_data[381]), .B0(n5587), .B1(
        image_data[509]), .Y(n5369) );
  NAND4XL U4317 ( .A(n5368), .B(n5367), .C(n5366), .D(n5365), .Y(n5374) );
  AOI22XL U4318 ( .A0(n5572), .A1(image_data[333]), .B0(n5571), .B1(
        image_data[461]), .Y(n5367) );
  AOI22XL U4319 ( .A0(n5574), .A1(image_data[301]), .B0(n5573), .B1(
        image_data[429]), .Y(n5366) );
  AOI22XL U4320 ( .A0(n5576), .A1(image_data[365]), .B0(n5575), .B1(
        image_data[493]), .Y(n5365) );
  NAND4XL U4321 ( .A(n5350), .B(n5349), .C(n5348), .D(n5347), .Y(n5351) );
  AOI22XL U4322 ( .A0(n5584), .A1(image_data[94]), .B0(n5583), .B1(
        image_data[222]), .Y(n5349) );
  AOI22XL U4323 ( .A0(n5586), .A1(image_data[62]), .B0(n5585), .B1(
        image_data[190]), .Y(n5348) );
  AOI22XL U4324 ( .A0(n5588), .A1(image_data[126]), .B0(n5587), .B1(
        image_data[254]), .Y(n5347) );
  NAND4XL U4325 ( .A(n5346), .B(n5345), .C(n5344), .D(n5343), .Y(n5352) );
  AOI22XL U4326 ( .A0(n5572), .A1(image_data[78]), .B0(n5571), .B1(
        image_data[206]), .Y(n5345) );
  AOI22XL U4327 ( .A0(n5574), .A1(image_data[46]), .B0(n5573), .B1(
        image_data[174]), .Y(n5344) );
  AOI22XL U4328 ( .A0(n5576), .A1(image_data[110]), .B0(n5575), .B1(
        image_data[238]), .Y(n5343) );
  NAND4XL U4329 ( .A(n5342), .B(n5341), .C(n5340), .D(n5339), .Y(n5353) );
  AOI22XL U4330 ( .A0(n5560), .A1(image_data[86]), .B0(n5559), .B1(
        image_data[214]), .Y(n5341) );
  AOI22XL U4331 ( .A0(n5562), .A1(image_data[54]), .B0(n5561), .B1(
        image_data[182]), .Y(n5340) );
  AOI22XL U4332 ( .A0(n5564), .A1(image_data[118]), .B0(n5563), .B1(
        image_data[246]), .Y(n5339) );
  NAND4XL U4333 ( .A(n5330), .B(n5329), .C(n5328), .D(n5327), .Y(n5331) );
  AOI22XL U4334 ( .A0(n5584), .A1(image_data[350]), .B0(n5583), .B1(
        image_data[478]), .Y(n5329) );
  AOI22XL U4335 ( .A0(n5586), .A1(image_data[318]), .B0(n5585), .B1(
        image_data[446]), .Y(n5328) );
  AOI22XL U4336 ( .A0(n5588), .A1(image_data[382]), .B0(n5587), .B1(
        image_data[510]), .Y(n5327) );
  NAND4XL U4337 ( .A(n5326), .B(n5325), .C(n5324), .D(n5323), .Y(n5332) );
  AOI22XL U4338 ( .A0(n5572), .A1(image_data[334]), .B0(n5571), .B1(
        image_data[462]), .Y(n5325) );
  AOI22XL U4339 ( .A0(n5574), .A1(image_data[302]), .B0(n5573), .B1(
        image_data[430]), .Y(n5324) );
  AOI22XL U4340 ( .A0(n5576), .A1(image_data[366]), .B0(n5575), .B1(
        image_data[494]), .Y(n5323) );
  NAND4XL U4341 ( .A(n5308), .B(n5307), .C(n5306), .D(n5305), .Y(n5309) );
  AOI22XL U4342 ( .A0(n5584), .A1(image_data[95]), .B0(n5583), .B1(
        image_data[223]), .Y(n5307) );
  AOI22XL U4343 ( .A0(n5586), .A1(image_data[63]), .B0(n5585), .B1(
        image_data[191]), .Y(n5306) );
  AOI22XL U4344 ( .A0(n5588), .A1(image_data[127]), .B0(n5587), .B1(
        image_data[255]), .Y(n5305) );
  NAND4XL U4345 ( .A(n5304), .B(n5303), .C(n5302), .D(n5301), .Y(n5310) );
  AOI22XL U4346 ( .A0(n5572), .A1(image_data[79]), .B0(n5571), .B1(
        image_data[207]), .Y(n5303) );
  AOI22XL U4347 ( .A0(n5574), .A1(image_data[47]), .B0(n5573), .B1(
        image_data[175]), .Y(n5302) );
  AOI22XL U4348 ( .A0(n5576), .A1(image_data[111]), .B0(n5575), .B1(
        image_data[239]), .Y(n5301) );
  NAND4XL U4349 ( .A(n5300), .B(n5299), .C(n5298), .D(n5297), .Y(n5311) );
  AOI22XL U4350 ( .A0(n5560), .A1(image_data[87]), .B0(n5559), .B1(
        image_data[215]), .Y(n5299) );
  AOI22XL U4351 ( .A0(n5562), .A1(image_data[55]), .B0(n5561), .B1(
        image_data[183]), .Y(n5298) );
  AOI22XL U4352 ( .A0(n5564), .A1(image_data[119]), .B0(n5563), .B1(
        image_data[247]), .Y(n5297) );
  NAND4XL U4353 ( .A(n5288), .B(n5287), .C(n5286), .D(n5285), .Y(n5289) );
  AOI22XL U4354 ( .A0(n5584), .A1(image_data[351]), .B0(n5583), .B1(
        image_data[479]), .Y(n5287) );
  AOI22XL U4355 ( .A0(n5586), .A1(image_data[319]), .B0(n5585), .B1(
        image_data[447]), .Y(n5286) );
  AOI22XL U4356 ( .A0(n5588), .A1(image_data[383]), .B0(n5587), .B1(
        image_data[511]), .Y(n5285) );
  NAND4XL U4357 ( .A(n5284), .B(n5283), .C(n5282), .D(n5281), .Y(n5290) );
  AOI22XL U4358 ( .A0(n5572), .A1(image_data[335]), .B0(n5571), .B1(
        image_data[463]), .Y(n5283) );
  AOI22XL U4359 ( .A0(n5574), .A1(image_data[303]), .B0(n5573), .B1(
        image_data[431]), .Y(n5282) );
  AOI22XL U4360 ( .A0(n5576), .A1(image_data[367]), .B0(n5575), .B1(
        image_data[495]), .Y(n5281) );
  OAI221XL U4361 ( .A0(in_valid), .A1(IRAM_D[0]), .B0(n8523), .B1(IROM_Q[0]), 
        .C0(n8480), .Y(n6121) );
  AOI22XL U4362 ( .A0(n6498), .A1(n6218), .B0(n6217), .B1(n6495), .Y(n6264) );
  OAI221XL U4363 ( .A0(in_valid), .A1(IRAM_D[1]), .B0(n8523), .B1(IROM_Q[1]), 
        .C0(n8480), .Y(n5696) );
  OAI21XL U4364 ( .A0(n6584), .A1(n6583), .B0(n6582), .Y(n6585) );
  AOI22XL U4365 ( .A0(n6498), .A1(n5082), .B0(n5081), .B1(n6495), .Y(n5265) );
  AOI222X1 U4366 ( .A0(n6581), .A1(n6018), .B0(n6579), .B1(n6017), .C0(n6577), 
        .C1(n6016), .Y(n6020) );
  CLKINVX3 U4367 ( .A(n8438), .Y(n8323) );
  NOR2X2 U4368 ( .A(n5185), .B(n5182), .Y(n5175) );
  NAND2XL U4369 ( .A(n4871), .B(n4985), .Y(n5097) );
  NOR2XL U4370 ( .A(n4871), .B(n4985), .Y(n5099) );
  INVXL U4371 ( .A(n8568), .Y(n4984) );
  NAND2XL U4372 ( .A(n5002), .B(n4588), .Y(n5171) );
  NOR2X2 U4373 ( .A(n5015), .B(n5012), .Y(n5005) );
  INVXL U4374 ( .A(n5178), .Y(n5180) );
  AOI2BB2XL U4375 ( .B0(op4[4]), .B1(n6131), .A0N(n6131), .A1N(op4[4]), .Y(
        n5184) );
  NOR2XL U4376 ( .A(N2760), .B(n4966), .Y(n5083) );
  NAND2BXL U4377 ( .AN(n4871), .B(n8458), .Y(n5084) );
  AOI22XL U4378 ( .A0(n8569), .A1(n4966), .B0(n8568), .B1(n4967), .Y(n5100) );
  NOR2XL U4379 ( .A(n8569), .B(n4966), .Y(n5102) );
  NAND2XL U4380 ( .A(n4871), .B(n5604), .Y(n5110) );
  INVXL U4381 ( .A(N2781), .Y(n4981) );
  INVXL U4382 ( .A(N2783), .Y(n4979) );
  NAND2XL U4383 ( .A(n8458), .B(n4985), .Y(n5135) );
  NOR2XL U4384 ( .A(n8458), .B(n4985), .Y(n5136) );
  AOI22XL U4385 ( .A0(n8569), .A1(n4986), .B0(n8568), .B1(n6173), .Y(n5137) );
  NOR2XL U4386 ( .A(n8569), .B(n4986), .Y(n5139) );
  INVXL U4387 ( .A(N2757), .Y(n4992) );
  INVX1 U4388 ( .A(N2779), .Y(n4978) );
  AOI22XL U4389 ( .A0(n6401), .A1(n5183), .B0(n5187), .B1(n8524), .Y(n5176) );
  INVX1 U4390 ( .A(n5195), .Y(n5191) );
  NOR2XL U4391 ( .A(N2774), .B(n5705), .Y(n5089) );
  AOI211XL U4392 ( .A0(n5088), .A1(n5087), .B0(n5086), .C0(n5085), .Y(n5090)
         );
  NAND2XL U4393 ( .A(N2779), .B(n5118), .Y(n5119) );
  AOI22XL U4394 ( .A0(n8567), .A1(n5115), .B0(n3442), .B1(n5118), .Y(n5106) );
  INVX1 U4395 ( .A(n5022), .Y(n5020) );
  INVX1 U4396 ( .A(n5023), .Y(n5019) );
  NAND2XL U4397 ( .A(n3470), .B(n8518), .Y(n3481) );
  AOI22XL U4398 ( .A0(n6550), .A1(image_data[104]), .B0(n6549), .B1(
        image_data[232]), .Y(n6102) );
  AOI22XL U4399 ( .A0(n6550), .A1(image_data[360]), .B0(n6549), .B1(
        image_data[488]), .Y(n6082) );
  AOI22XL U4400 ( .A0(n6474), .A1(image_data[104]), .B0(n6473), .B1(
        image_data[232]), .Y(n6060) );
  AOI22XL U4401 ( .A0(n6550), .A1(image_data[110]), .B0(n6549), .B1(
        image_data[238]), .Y(n5883) );
  AOI22XL U4402 ( .A0(n6550), .A1(image_data[366]), .B0(n6549), .B1(
        image_data[494]), .Y(n5863) );
  AOI22XL U4403 ( .A0(n6474), .A1(image_data[110]), .B0(n6473), .B1(
        image_data[238]), .Y(n5841) );
  AOI22XL U4404 ( .A0(n6550), .A1(image_data[105]), .B0(n6549), .B1(
        image_data[233]), .Y(n5678) );
  AOI22XL U4405 ( .A0(n6550), .A1(image_data[361]), .B0(n6549), .B1(
        image_data[489]), .Y(n5658) );
  AOI22XL U4406 ( .A0(n6474), .A1(image_data[105]), .B0(n6473), .B1(
        image_data[233]), .Y(n5636) );
  AOI22XL U4407 ( .A0(n6550), .A1(image_data[108]), .B0(n6549), .B1(
        image_data[236]), .Y(n5780) );
  AOI22XL U4408 ( .A0(n6550), .A1(image_data[364]), .B0(n6549), .B1(
        image_data[492]), .Y(n5760) );
  AOI22XL U4409 ( .A0(n6474), .A1(image_data[108]), .B0(n6473), .B1(
        image_data[236]), .Y(n5738) );
  NOR2XL U4410 ( .A(n8569), .B(n4872), .Y(n4780) );
  NOR2XL U4411 ( .A(n3442), .B(n4978), .Y(n5162) );
  NAND2XL U4412 ( .A(N2755), .B(n4978), .Y(n5149) );
  NAND2XL U4413 ( .A(N2755), .B(n3441), .Y(n5148) );
  AOI22XL U4414 ( .A0(n3895), .A1(image_data[66]), .B0(n3364), .B1(
        image_data[194]), .Y(n3795) );
  AOI22XL U4415 ( .A0(n3878), .A1(image_data[122]), .B0(n3811), .B1(
        image_data[250]), .Y(n3812) );
  AOI22XL U4416 ( .A0(n3868), .A1(image_data[106]), .B0(n3805), .B1(
        image_data[234]), .Y(n3806) );
  AOI22XL U4417 ( .A0(n3935), .A1(image_data[114]), .B0(n3799), .B1(
        image_data[242]), .Y(n3800) );
  AOI22XL U4418 ( .A0(n3895), .A1(image_data[322]), .B0(n3364), .B1(
        image_data[450]), .Y(n3773) );
  AOI22XL U4419 ( .A0(n3878), .A1(image_data[378]), .B0(n3879), .B1(
        image_data[506]), .Y(n3783) );
  AOI22XL U4420 ( .A0(n3868), .A1(image_data[362]), .B0(n3869), .B1(
        image_data[490]), .Y(n3779) );
  NAND2XL U4421 ( .A(n5215), .B(n5214), .Y(n5223) );
  NAND2XL U4422 ( .A(n5215), .B(n5208), .Y(n5209) );
  NAND2XL U4423 ( .A(n5202), .B(n5208), .Y(n5197) );
  OAI21XL U4424 ( .A0(n5108), .A1(n5107), .B0(n5106), .Y(n5123) );
  OAI21XL U4425 ( .A0(n5121), .A1(n5120), .B0(n5119), .Y(n5122) );
  AOI22XL U4426 ( .A0(n5096), .A1(n5095), .B0(N2755), .B1(n5118), .Y(n5125) );
  OAI21XL U4427 ( .A0(n5162), .A1(n5161), .B0(n5160), .Y(n5163) );
  AOI22XL U4428 ( .A0(n5159), .A1(n5158), .B0(n8567), .B1(n5807), .Y(n5161) );
  AOI21XL U4429 ( .A0(n5154), .A1(n5153), .B0(n5152), .Y(n5157) );
  AOI21XL U4430 ( .A0(n5142), .A1(n5141), .B0(n5140), .Y(n5145) );
  NAND2XL U4431 ( .A(n5043), .B(n5042), .Y(n5051) );
  NAND2XL U4432 ( .A(n5043), .B(n5036), .Y(n5037) );
  NAND2XL U4433 ( .A(n5030), .B(n5036), .Y(n5025) );
  NAND3XL U4434 ( .A(op4[4]), .B(op2[2]), .C(n6401), .Y(n3487) );
  AOI22XL U4435 ( .A0(n3364), .A1(image_data[0]), .B0(n3895), .B1(
        image_data[128]), .Y(n4619) );
  NAND3XL U4436 ( .A(op4[4]), .B(n6401), .C(n8528), .Y(n3484) );
  AOI22XL U4437 ( .A0(n3878), .A1(image_data[123]), .B0(n3811), .B1(
        image_data[251]), .Y(n3761) );
  AOI22XL U4438 ( .A0(n3893), .A1(image_data[99]), .B0(n3792), .B1(
        image_data[227]), .Y(n3749) );
  AOI22XL U4439 ( .A0(n3868), .A1(image_data[107]), .B0(n3805), .B1(
        image_data[235]), .Y(n3757) );
  NOR2X1 U4440 ( .A(n3486), .B(n3471), .Y(n3798) );
  AOI22XL U4441 ( .A0(n3935), .A1(image_data[115]), .B0(n3799), .B1(
        image_data[243]), .Y(n3753) );
  AOI22XL U4442 ( .A0(n3878), .A1(image_data[379]), .B0(n3811), .B1(
        image_data[507]), .Y(n3741) );
  AOI22XL U4443 ( .A0(n3893), .A1(image_data[355]), .B0(n3792), .B1(
        image_data[483]), .Y(n3729) );
  AOI22XL U4444 ( .A0(n3868), .A1(image_data[363]), .B0(n3805), .B1(
        image_data[491]), .Y(n3737) );
  AOI22XL U4445 ( .A0(n3874), .A1(image_data[95]), .B0(n3948), .B1(
        image_data[223]), .Y(n3510) );
  AOI22XL U4446 ( .A0(n3942), .A1(image_data[111]), .B0(n3943), .B1(
        image_data[239]), .Y(n3504) );
  AOI22XL U4447 ( .A0(n3884), .A1(image_data[87]), .B0(n3934), .B1(
        image_data[215]), .Y(n3502) );
  AOI22XL U4448 ( .A0(n3894), .A1(image_data[39]), .B0(n3893), .B1(
        image_data[167]), .Y(n3497) );
  AOI22XL U4449 ( .A0(n3874), .A1(image_data[351]), .B0(n3948), .B1(
        image_data[479]), .Y(n3490) );
  AOI22XL U4450 ( .A0(n4754), .A1(image_data[367]), .B0(n3943), .B1(
        image_data[495]), .Y(n3477) );
  AOI22XL U4451 ( .A0(n3884), .A1(image_data[343]), .B0(n3934), .B1(
        image_data[471]), .Y(n3474) );
  AOI22XL U4452 ( .A0(n3894), .A1(image_data[295]), .B0(n3893), .B1(
        image_data[423]), .Y(n3467) );
  AND3XL U4453 ( .A(op2[2]), .B(op4[4]), .C(n8524), .Y(n3401) );
  AND2XL U4454 ( .A(IROM_A[0]), .B(n8520), .Y(n3402) );
  AND2XL U4455 ( .A(IROM_A[1]), .B(n8526), .Y(n3403) );
  AOI22XL U4456 ( .A0(n3895), .A1(image_data[65]), .B0(n3364), .B1(
        image_data[193]), .Y(n4941) );
  AOI22XL U4457 ( .A0(n3874), .A1(image_data[25]), .B0(n3948), .B1(
        image_data[153]), .Y(n4954) );
  AOI22XL U4458 ( .A0(n3887), .A1(image_data[49]), .B0(n3936), .B1(
        image_data[177]), .Y(n4944) );
  AOI22XL U4459 ( .A0(n3942), .A1(image_data[41]), .B0(n3943), .B1(
        image_data[169]), .Y(n4948) );
  AOI22XL U4460 ( .A0(n3895), .A1(image_data[321]), .B0(n3364), .B1(
        image_data[449]), .Y(n4921) );
  AOI22XL U4461 ( .A0(n3878), .A1(image_data[377]), .B0(n3879), .B1(
        image_data[505]), .Y(n4931) );
  AOI22XL U4462 ( .A0(n3868), .A1(image_data[361]), .B0(n3869), .B1(
        image_data[489]), .Y(n4927) );
  AOI22XL U4463 ( .A0(n3895), .A1(image_data[121]), .B0(n3364), .B1(
        image_data[249]), .Y(n4671) );
  AOI22XL U4464 ( .A0(n3879), .A1(image_data[49]), .B0(n3878), .B1(
        image_data[177]), .Y(n4663) );
  AOI22XL U4465 ( .A0(n3869), .A1(image_data[33]), .B0(n3868), .B1(
        image_data[161]), .Y(n4659) );
  AOI22XL U4466 ( .A0(n3884), .A1(image_data[73]), .B0(n3934), .B1(
        image_data[201]), .Y(n4668) );
  AOI22XL U4467 ( .A0(n3895), .A1(image_data[377]), .B0(n3364), .B1(
        image_data[505]), .Y(n4650) );
  AOI22XL U4468 ( .A0(n3879), .A1(image_data[305]), .B0(n3878), .B1(
        image_data[433]), .Y(n4643) );
  AOI22XL U4469 ( .A0(n3869), .A1(image_data[289]), .B0(n3868), .B1(
        image_data[417]), .Y(n4639) );
  AOI22XL U4470 ( .A0(n3935), .A1(image_data[112]), .B0(n3888), .B1(
        image_data[240]), .Y(n4901) );
  AOI22XL U4471 ( .A0(n3895), .A1(image_data[64]), .B0(n3364), .B1(
        image_data[192]), .Y(n4899) );
  AOI22XL U4472 ( .A0(n4714), .A1(image_data[104]), .B0(n3869), .B1(
        image_data[232]), .Y(n4905) );
  AOI22XL U4473 ( .A0(n4721), .A1(image_data[120]), .B0(n3879), .B1(
        image_data[248]), .Y(n4909) );
  AOI22XL U4474 ( .A0(n3935), .A1(image_data[368]), .B0(n3888), .B1(
        image_data[496]), .Y(n4881) );
  AOI22XL U4475 ( .A0(n3895), .A1(image_data[320]), .B0(n3364), .B1(
        image_data[448]), .Y(n4879) );
  AOI22XL U4476 ( .A0(n4714), .A1(image_data[360]), .B0(n3869), .B1(
        image_data[488]), .Y(n4885) );
  AOI22XL U4477 ( .A0(n3895), .A1(image_data[120]), .B0(n3364), .B1(
        image_data[248]), .Y(n4769) );
  AOI22XL U4478 ( .A0(n3879), .A1(image_data[48]), .B0(n3878), .B1(
        image_data[176]), .Y(n4760) );
  AOI22XL U4479 ( .A0(n3869), .A1(image_data[32]), .B0(n3868), .B1(
        image_data[160]), .Y(n4756) );
  AOI22XL U4480 ( .A0(n3884), .A1(image_data[72]), .B0(n3934), .B1(
        image_data[200]), .Y(n4766) );
  AOI22XL U4481 ( .A0(n3879), .A1(image_data[304]), .B0(n3878), .B1(
        image_data[432]), .Y(n4738) );
  AOI22XL U4482 ( .A0(n3894), .A1(image_data[280]), .B0(n3893), .B1(
        image_data[408]), .Y(n4748) );
  AOI22XL U4483 ( .A0(n3869), .A1(image_data[288]), .B0(n3868), .B1(
        image_data[416]), .Y(n4734) );
  OAI2BB1XL U4484 ( .A0N(n6124), .A1N(n5258), .B0(n5257), .Y(n5261) );
  AOI22XL U4485 ( .A0(n6474), .A1(image_data[360]), .B0(n6473), .B1(
        image_data[488]), .Y(n6040) );
  AOI22XL U4486 ( .A0(n6486), .A1(image_data[376]), .B0(n6485), .B1(
        image_data[504]), .Y(n6044) );
  AOI22XL U4487 ( .A0(n6450), .A1(image_data[352]), .B0(n6449), .B1(
        image_data[480]), .Y(n6032) );
  AOI22XL U4488 ( .A0(n6458), .A1(image_data[336]), .B0(n6457), .B1(
        image_data[464]), .Y(n6038) );
  AOI22XL U4489 ( .A0(n6562), .A1(image_data[120]), .B0(n6561), .B1(
        image_data[248]), .Y(n6106) );
  AOI22XL U4490 ( .A0(n6560), .A1(image_data[56]), .B0(n6559), .B1(
        image_data[184]), .Y(n6107) );
  AOI22XL U4491 ( .A0(n6558), .A1(image_data[88]), .B0(n6557), .B1(
        image_data[216]), .Y(n6108) );
  AOI22XL U4492 ( .A0(n6556), .A1(image_data[24]), .B0(n6555), .B1(
        image_data[152]), .Y(n6109) );
  AOI22XL U4493 ( .A0(n6526), .A1(image_data[96]), .B0(n6525), .B1(
        image_data[224]), .Y(n6094) );
  AOI22XL U4494 ( .A0(n6524), .A1(image_data[32]), .B0(n6523), .B1(
        image_data[160]), .Y(n6095) );
  AOI22XL U4495 ( .A0(n6522), .A1(image_data[64]), .B0(n6521), .B1(
        image_data[192]), .Y(n6096) );
  AOI22XL U4496 ( .A0(n6520), .A1(image_data[0]), .B0(n6519), .B1(
        image_data[128]), .Y(n6097) );
  AOI22XL U4497 ( .A0(n6534), .A1(image_data[80]), .B0(n6533), .B1(
        image_data[208]), .Y(n6100) );
  AOI22XL U4498 ( .A0(n6538), .A1(image_data[112]), .B0(n6537), .B1(
        image_data[240]), .Y(n6098) );
  AOI22XL U4499 ( .A0(n6536), .A1(image_data[48]), .B0(n6535), .B1(
        image_data[176]), .Y(n6099) );
  AOI22XL U4500 ( .A0(n6532), .A1(image_data[16]), .B0(n6531), .B1(
        image_data[144]), .Y(n6101) );
  NAND4XL U4501 ( .A(n6105), .B(n6104), .C(n6103), .D(n6102), .Y(n6111) );
  AOI22XL U4502 ( .A0(n6544), .A1(image_data[8]), .B0(n6543), .B1(
        image_data[136]), .Y(n6105) );
  AOI22XL U4503 ( .A0(n6546), .A1(image_data[72]), .B0(n6545), .B1(
        image_data[200]), .Y(n6104) );
  AOI22XL U4504 ( .A0(n6548), .A1(image_data[40]), .B0(n6547), .B1(
        image_data[168]), .Y(n6103) );
  AOI22XL U4505 ( .A0(n6562), .A1(image_data[376]), .B0(n6561), .B1(
        image_data[504]), .Y(n6086) );
  AOI22XL U4506 ( .A0(n6560), .A1(image_data[312]), .B0(n6559), .B1(
        image_data[440]), .Y(n6087) );
  AOI22XL U4507 ( .A0(n6558), .A1(image_data[344]), .B0(n6557), .B1(
        image_data[472]), .Y(n6088) );
  AOI22XL U4508 ( .A0(n6556), .A1(image_data[280]), .B0(n6555), .B1(
        image_data[408]), .Y(n6089) );
  AOI22XL U4509 ( .A0(n6526), .A1(image_data[352]), .B0(n6525), .B1(
        image_data[480]), .Y(n6074) );
  AOI22XL U4510 ( .A0(n6524), .A1(image_data[288]), .B0(n6523), .B1(
        image_data[416]), .Y(n6075) );
  AOI22XL U4511 ( .A0(n6522), .A1(image_data[320]), .B0(n6521), .B1(
        image_data[448]), .Y(n6076) );
  AOI22XL U4512 ( .A0(n6520), .A1(image_data[256]), .B0(n6519), .B1(
        image_data[384]), .Y(n6077) );
  AOI22XL U4513 ( .A0(n6534), .A1(image_data[336]), .B0(n6533), .B1(
        image_data[464]), .Y(n6080) );
  AOI22XL U4514 ( .A0(n6538), .A1(image_data[368]), .B0(n6537), .B1(
        image_data[496]), .Y(n6078) );
  AOI22XL U4515 ( .A0(n6536), .A1(image_data[304]), .B0(n6535), .B1(
        image_data[432]), .Y(n6079) );
  AOI22XL U4516 ( .A0(n6532), .A1(image_data[272]), .B0(n6531), .B1(
        image_data[400]), .Y(n6081) );
  NAND4XL U4517 ( .A(n6085), .B(n6084), .C(n6083), .D(n6082), .Y(n6091) );
  AOI22XL U4518 ( .A0(n6544), .A1(image_data[264]), .B0(n6543), .B1(
        image_data[392]), .Y(n6085) );
  AOI22XL U4519 ( .A0(n6546), .A1(image_data[328]), .B0(n6545), .B1(
        image_data[456]), .Y(n6084) );
  AOI22XL U4520 ( .A0(n6548), .A1(image_data[296]), .B0(n6547), .B1(
        image_data[424]), .Y(n6083) );
  AOI22XL U4521 ( .A0(n6486), .A1(image_data[120]), .B0(n6485), .B1(
        image_data[248]), .Y(n6064) );
  AOI22XL U4522 ( .A0(n6484), .A1(image_data[56]), .B0(n6483), .B1(
        image_data[184]), .Y(n6065) );
  AOI22XL U4523 ( .A0(n6482), .A1(image_data[88]), .B0(n6481), .B1(
        image_data[216]), .Y(n6066) );
  AOI22XL U4524 ( .A0(n6480), .A1(image_data[24]), .B0(n6479), .B1(
        image_data[152]), .Y(n6067) );
  AOI22XL U4525 ( .A0(n6450), .A1(image_data[96]), .B0(n6449), .B1(
        image_data[224]), .Y(n6052) );
  AOI22XL U4526 ( .A0(n6448), .A1(image_data[32]), .B0(n6447), .B1(
        image_data[160]), .Y(n6053) );
  AOI22XL U4527 ( .A0(n6446), .A1(image_data[64]), .B0(n6445), .B1(
        image_data[192]), .Y(n6054) );
  AOI22XL U4528 ( .A0(n6444), .A1(image_data[0]), .B0(n6443), .B1(
        image_data[128]), .Y(n6055) );
  AOI22XL U4529 ( .A0(n6458), .A1(image_data[80]), .B0(n6457), .B1(
        image_data[208]), .Y(n6058) );
  AOI22XL U4530 ( .A0(n6462), .A1(image_data[112]), .B0(n6461), .B1(
        image_data[240]), .Y(n6056) );
  AOI22XL U4531 ( .A0(n6460), .A1(image_data[48]), .B0(n6459), .B1(
        image_data[176]), .Y(n6057) );
  AOI22XL U4532 ( .A0(n6456), .A1(image_data[16]), .B0(n6455), .B1(
        image_data[144]), .Y(n6059) );
  NAND4XL U4533 ( .A(n6063), .B(n6062), .C(n6061), .D(n6060), .Y(n6069) );
  AOI22XL U4534 ( .A0(n6468), .A1(image_data[8]), .B0(n6467), .B1(
        image_data[136]), .Y(n6063) );
  AOI22XL U4535 ( .A0(n6470), .A1(image_data[72]), .B0(n6469), .B1(
        image_data[200]), .Y(n6062) );
  AOI22XL U4536 ( .A0(n6472), .A1(image_data[40]), .B0(n6471), .B1(
        image_data[168]), .Y(n6061) );
  AOI22XL U4537 ( .A0(n3895), .A1(image_data[57]), .B0(n3364), .B1(
        image_data[185]), .Y(n4861) );
  AOI22XL U4538 ( .A0(n3887), .A1(image_data[41]), .B0(n3936), .B1(
        image_data[169]), .Y(n4857) );
  AOI22XL U4539 ( .A0(n3878), .A1(image_data[113]), .B0(n3879), .B1(
        image_data[241]), .Y(n4852) );
  AOI22XL U4540 ( .A0(n3868), .A1(image_data[97]), .B0(n3869), .B1(
        image_data[225]), .Y(n4848) );
  AOI22XL U4541 ( .A0(n3895), .A1(image_data[313]), .B0(n3364), .B1(
        image_data[441]), .Y(n4841) );
  AOI22XL U4542 ( .A0(n3887), .A1(image_data[297]), .B0(n3936), .B1(
        image_data[425]), .Y(n4837) );
  AOI22XL U4543 ( .A0(n3878), .A1(image_data[369]), .B0(n3879), .B1(
        image_data[497]), .Y(n4832) );
  AOI22XL U4544 ( .A0(n3868), .A1(image_data[353]), .B0(n3869), .B1(
        image_data[481]), .Y(n4828) );
  AOI22XL U4545 ( .A0(n3364), .A1(image_data[1]), .B0(n3895), .B1(
        image_data[129]), .Y(n4706) );
  AOI22XL U4546 ( .A0(n4720), .A1(image_data[89]), .B0(n3948), .B1(
        image_data[217]), .Y(n4725) );
  AOI22XL U4547 ( .A0(n3942), .A1(image_data[105]), .B0(n3943), .B1(
        image_data[233]), .Y(n4715) );
  AOI22XL U4548 ( .A0(n4708), .A1(image_data[81]), .B0(n3934), .B1(
        image_data[209]), .Y(n4711) );
  AOI22XL U4549 ( .A0(n4720), .A1(image_data[345]), .B0(n3948), .B1(
        image_data[473]), .Y(n4696) );
  AOI22XL U4550 ( .A0(n3942), .A1(image_data[361]), .B0(n3943), .B1(
        image_data[489]), .Y(n4690) );
  AOI22XL U4551 ( .A0(n3894), .A1(image_data[289]), .B0(n3893), .B1(
        image_data[417]), .Y(n4683) );
  AOI22XL U4552 ( .A0(n6474), .A1(image_data[107]), .B0(n6473), .B1(
        image_data[235]), .Y(n6205) );
  AOI22XL U4553 ( .A0(n6474), .A1(image_data[363]), .B0(n6473), .B1(
        image_data[491]), .Y(n6185) );
  AOI22XL U4554 ( .A0(n6550), .A1(image_data[107]), .B0(n6549), .B1(
        image_data[235]), .Y(n6247) );
  AOI22XL U4555 ( .A0(n6562), .A1(image_data[123]), .B0(n6561), .B1(
        image_data[251]), .Y(n6251) );
  AOI22XL U4556 ( .A0(n6526), .A1(image_data[99]), .B0(n6525), .B1(
        image_data[227]), .Y(n6239) );
  AOI22XL U4557 ( .A0(n6534), .A1(image_data[83]), .B0(n6533), .B1(
        image_data[211]), .Y(n6245) );
  AOI22XL U4558 ( .A0(n6550), .A1(image_data[363]), .B0(n6549), .B1(
        image_data[491]), .Y(n6227) );
  AOI22XL U4559 ( .A0(n6562), .A1(image_data[379]), .B0(n6561), .B1(
        image_data[507]), .Y(n6231) );
  AOI22XL U4560 ( .A0(n6526), .A1(image_data[355]), .B0(n6525), .B1(
        image_data[483]), .Y(n6219) );
  AOI22XL U4561 ( .A0(n6474), .A1(image_data[366]), .B0(n6473), .B1(
        image_data[494]), .Y(n5821) );
  AOI22XL U4562 ( .A0(n6486), .A1(image_data[382]), .B0(n6485), .B1(
        image_data[510]), .Y(n5825) );
  AOI22XL U4563 ( .A0(n6450), .A1(image_data[358]), .B0(n6449), .B1(
        image_data[486]), .Y(n5813) );
  AOI22XL U4564 ( .A0(n6458), .A1(image_data[342]), .B0(n6457), .B1(
        image_data[470]), .Y(n5819) );
  AOI22XL U4565 ( .A0(n6562), .A1(image_data[126]), .B0(n6561), .B1(
        image_data[254]), .Y(n5887) );
  AOI22XL U4566 ( .A0(n6560), .A1(image_data[62]), .B0(n6559), .B1(
        image_data[190]), .Y(n5888) );
  AOI22XL U4567 ( .A0(n6558), .A1(image_data[94]), .B0(n6557), .B1(
        image_data[222]), .Y(n5889) );
  AOI22XL U4568 ( .A0(n6556), .A1(image_data[30]), .B0(n6555), .B1(
        image_data[158]), .Y(n5890) );
  AOI22XL U4569 ( .A0(n6526), .A1(image_data[102]), .B0(n6525), .B1(
        image_data[230]), .Y(n5875) );
  AOI22XL U4570 ( .A0(n6524), .A1(image_data[38]), .B0(n6523), .B1(
        image_data[166]), .Y(n5876) );
  AOI22XL U4571 ( .A0(n6522), .A1(image_data[70]), .B0(n6521), .B1(
        image_data[198]), .Y(n5877) );
  AOI22XL U4572 ( .A0(n6520), .A1(image_data[6]), .B0(n6519), .B1(
        image_data[134]), .Y(n5878) );
  AOI22XL U4573 ( .A0(n6534), .A1(image_data[86]), .B0(n6533), .B1(
        image_data[214]), .Y(n5881) );
  AOI22XL U4574 ( .A0(n6538), .A1(image_data[118]), .B0(n6537), .B1(
        image_data[246]), .Y(n5879) );
  AOI22XL U4575 ( .A0(n6536), .A1(image_data[54]), .B0(n6535), .B1(
        image_data[182]), .Y(n5880) );
  AOI22XL U4576 ( .A0(n6532), .A1(image_data[22]), .B0(n6531), .B1(
        image_data[150]), .Y(n5882) );
  NAND4XL U4577 ( .A(n5886), .B(n5885), .C(n5884), .D(n5883), .Y(n5892) );
  AOI22XL U4578 ( .A0(n6544), .A1(image_data[14]), .B0(n6543), .B1(
        image_data[142]), .Y(n5886) );
  AOI22XL U4579 ( .A0(n6546), .A1(image_data[78]), .B0(n6545), .B1(
        image_data[206]), .Y(n5885) );
  AOI22XL U4580 ( .A0(n6548), .A1(image_data[46]), .B0(n6547), .B1(
        image_data[174]), .Y(n5884) );
  AOI22XL U4581 ( .A0(n6562), .A1(image_data[382]), .B0(n6561), .B1(
        image_data[510]), .Y(n5867) );
  AOI22XL U4582 ( .A0(n6560), .A1(image_data[318]), .B0(n6559), .B1(
        image_data[446]), .Y(n5868) );
  AOI22XL U4583 ( .A0(n6558), .A1(image_data[350]), .B0(n6557), .B1(
        image_data[478]), .Y(n5869) );
  AOI22XL U4584 ( .A0(n6556), .A1(image_data[286]), .B0(n6555), .B1(
        image_data[414]), .Y(n5870) );
  AOI22XL U4585 ( .A0(n6526), .A1(image_data[358]), .B0(n6525), .B1(
        image_data[486]), .Y(n5855) );
  AOI22XL U4586 ( .A0(n6524), .A1(image_data[294]), .B0(n6523), .B1(
        image_data[422]), .Y(n5856) );
  AOI22XL U4587 ( .A0(n6522), .A1(image_data[326]), .B0(n6521), .B1(
        image_data[454]), .Y(n5857) );
  AOI22XL U4588 ( .A0(n6520), .A1(image_data[262]), .B0(n6519), .B1(
        image_data[390]), .Y(n5858) );
  AOI22XL U4589 ( .A0(n6534), .A1(image_data[342]), .B0(n6533), .B1(
        image_data[470]), .Y(n5861) );
  AOI22XL U4590 ( .A0(n6538), .A1(image_data[374]), .B0(n6537), .B1(
        image_data[502]), .Y(n5859) );
  AOI22XL U4591 ( .A0(n6536), .A1(image_data[310]), .B0(n6535), .B1(
        image_data[438]), .Y(n5860) );
  AOI22XL U4592 ( .A0(n6532), .A1(image_data[278]), .B0(n6531), .B1(
        image_data[406]), .Y(n5862) );
  NAND4XL U4593 ( .A(n5866), .B(n5865), .C(n5864), .D(n5863), .Y(n5872) );
  AOI22XL U4594 ( .A0(n6544), .A1(image_data[270]), .B0(n6543), .B1(
        image_data[398]), .Y(n5866) );
  AOI22XL U4595 ( .A0(n6546), .A1(image_data[334]), .B0(n6545), .B1(
        image_data[462]), .Y(n5865) );
  AOI22XL U4596 ( .A0(n6548), .A1(image_data[302]), .B0(n6547), .B1(
        image_data[430]), .Y(n5864) );
  AOI22XL U4597 ( .A0(n6486), .A1(image_data[126]), .B0(n6485), .B1(
        image_data[254]), .Y(n5845) );
  AOI22XL U4598 ( .A0(n6484), .A1(image_data[62]), .B0(n6483), .B1(
        image_data[190]), .Y(n5846) );
  AOI22XL U4599 ( .A0(n6482), .A1(image_data[94]), .B0(n6481), .B1(
        image_data[222]), .Y(n5847) );
  AOI22XL U4600 ( .A0(n6480), .A1(image_data[30]), .B0(n6479), .B1(
        image_data[158]), .Y(n5848) );
  AOI22XL U4601 ( .A0(n6450), .A1(image_data[102]), .B0(n6449), .B1(
        image_data[230]), .Y(n5833) );
  AOI22XL U4602 ( .A0(n6448), .A1(image_data[38]), .B0(n6447), .B1(
        image_data[166]), .Y(n5834) );
  AOI22XL U4603 ( .A0(n6446), .A1(image_data[70]), .B0(n6445), .B1(
        image_data[198]), .Y(n5835) );
  AOI22XL U4604 ( .A0(n6444), .A1(image_data[6]), .B0(n6443), .B1(
        image_data[134]), .Y(n5836) );
  AOI22XL U4605 ( .A0(n6458), .A1(image_data[86]), .B0(n6457), .B1(
        image_data[214]), .Y(n5839) );
  AOI22XL U4606 ( .A0(n6462), .A1(image_data[118]), .B0(n6461), .B1(
        image_data[246]), .Y(n5837) );
  AOI22XL U4607 ( .A0(n6460), .A1(image_data[54]), .B0(n6459), .B1(
        image_data[182]), .Y(n5838) );
  AOI22XL U4608 ( .A0(n6456), .A1(image_data[22]), .B0(n6455), .B1(
        image_data[150]), .Y(n5840) );
  NAND4XL U4609 ( .A(n5844), .B(n5843), .C(n5842), .D(n5841), .Y(n5850) );
  AOI22XL U4610 ( .A0(n6468), .A1(image_data[14]), .B0(n6467), .B1(
        image_data[142]), .Y(n5844) );
  AOI22XL U4611 ( .A0(n6470), .A1(image_data[78]), .B0(n6469), .B1(
        image_data[206]), .Y(n5843) );
  AOI22XL U4612 ( .A0(n6472), .A1(image_data[46]), .B0(n6471), .B1(
        image_data[174]), .Y(n5842) );
  AOI22XL U4613 ( .A0(n6474), .A1(image_data[361]), .B0(n6473), .B1(
        image_data[489]), .Y(n5616) );
  AOI22XL U4614 ( .A0(n6486), .A1(image_data[377]), .B0(n6485), .B1(
        image_data[505]), .Y(n5620) );
  AOI22XL U4615 ( .A0(n6450), .A1(image_data[353]), .B0(n6449), .B1(
        image_data[481]), .Y(n5608) );
  AOI22XL U4616 ( .A0(n6458), .A1(image_data[337]), .B0(n6457), .B1(
        image_data[465]), .Y(n5614) );
  AOI22XL U4617 ( .A0(n6562), .A1(image_data[121]), .B0(n6561), .B1(
        image_data[249]), .Y(n5682) );
  AOI22XL U4618 ( .A0(n6560), .A1(image_data[57]), .B0(n6559), .B1(
        image_data[185]), .Y(n5683) );
  AOI22XL U4619 ( .A0(n6558), .A1(image_data[89]), .B0(n6557), .B1(
        image_data[217]), .Y(n5684) );
  AOI22XL U4620 ( .A0(n6556), .A1(image_data[25]), .B0(n6555), .B1(
        image_data[153]), .Y(n5685) );
  AOI22XL U4621 ( .A0(n6526), .A1(image_data[97]), .B0(n6525), .B1(
        image_data[225]), .Y(n5670) );
  AOI22XL U4622 ( .A0(n6524), .A1(image_data[33]), .B0(n6523), .B1(
        image_data[161]), .Y(n5671) );
  AOI22XL U4623 ( .A0(n6522), .A1(image_data[65]), .B0(n6521), .B1(
        image_data[193]), .Y(n5672) );
  AOI22XL U4624 ( .A0(n6520), .A1(image_data[1]), .B0(n6519), .B1(
        image_data[129]), .Y(n5673) );
  AOI22XL U4625 ( .A0(n6534), .A1(image_data[81]), .B0(n6533), .B1(
        image_data[209]), .Y(n5676) );
  AOI22XL U4626 ( .A0(n6538), .A1(image_data[113]), .B0(n6537), .B1(
        image_data[241]), .Y(n5674) );
  AOI22XL U4627 ( .A0(n6536), .A1(image_data[49]), .B0(n6535), .B1(
        image_data[177]), .Y(n5675) );
  AOI22XL U4628 ( .A0(n6532), .A1(image_data[17]), .B0(n6531), .B1(
        image_data[145]), .Y(n5677) );
  NAND4XL U4629 ( .A(n5681), .B(n5680), .C(n5679), .D(n5678), .Y(n5687) );
  AOI22XL U4630 ( .A0(n6544), .A1(image_data[9]), .B0(n6543), .B1(
        image_data[137]), .Y(n5681) );
  AOI22XL U4631 ( .A0(n6546), .A1(image_data[73]), .B0(n6545), .B1(
        image_data[201]), .Y(n5680) );
  AOI22XL U4632 ( .A0(n6548), .A1(image_data[41]), .B0(n6547), .B1(
        image_data[169]), .Y(n5679) );
  AOI22XL U4633 ( .A0(n6562), .A1(image_data[377]), .B0(n6561), .B1(
        image_data[505]), .Y(n5662) );
  AOI22XL U4634 ( .A0(n6560), .A1(image_data[313]), .B0(n6559), .B1(
        image_data[441]), .Y(n5663) );
  AOI22XL U4635 ( .A0(n6558), .A1(image_data[345]), .B0(n6557), .B1(
        image_data[473]), .Y(n5664) );
  AOI22XL U4636 ( .A0(n6556), .A1(image_data[281]), .B0(n6555), .B1(
        image_data[409]), .Y(n5665) );
  AOI22XL U4637 ( .A0(n6526), .A1(image_data[353]), .B0(n6525), .B1(
        image_data[481]), .Y(n5650) );
  AOI22XL U4638 ( .A0(n6524), .A1(image_data[289]), .B0(n6523), .B1(
        image_data[417]), .Y(n5651) );
  AOI22XL U4639 ( .A0(n6522), .A1(image_data[321]), .B0(n6521), .B1(
        image_data[449]), .Y(n5652) );
  AOI22XL U4640 ( .A0(n6520), .A1(image_data[257]), .B0(n6519), .B1(
        image_data[385]), .Y(n5653) );
  AOI22XL U4641 ( .A0(n6534), .A1(image_data[337]), .B0(n6533), .B1(
        image_data[465]), .Y(n5656) );
  AOI22XL U4642 ( .A0(n6538), .A1(image_data[369]), .B0(n6537), .B1(
        image_data[497]), .Y(n5654) );
  AOI22XL U4643 ( .A0(n6536), .A1(image_data[305]), .B0(n6535), .B1(
        image_data[433]), .Y(n5655) );
  AOI22XL U4644 ( .A0(n6532), .A1(image_data[273]), .B0(n6531), .B1(
        image_data[401]), .Y(n5657) );
  NAND4XL U4645 ( .A(n5661), .B(n5660), .C(n5659), .D(n5658), .Y(n5667) );
  AOI22XL U4646 ( .A0(n6544), .A1(image_data[265]), .B0(n6543), .B1(
        image_data[393]), .Y(n5661) );
  AOI22XL U4647 ( .A0(n6546), .A1(image_data[329]), .B0(n6545), .B1(
        image_data[457]), .Y(n5660) );
  AOI22XL U4648 ( .A0(n6548), .A1(image_data[297]), .B0(n6547), .B1(
        image_data[425]), .Y(n5659) );
  AOI22XL U4649 ( .A0(n6486), .A1(image_data[121]), .B0(n6485), .B1(
        image_data[249]), .Y(n5640) );
  AOI22XL U4650 ( .A0(n6484), .A1(image_data[57]), .B0(n6483), .B1(
        image_data[185]), .Y(n5641) );
  AOI22XL U4651 ( .A0(n6482), .A1(image_data[89]), .B0(n6481), .B1(
        image_data[217]), .Y(n5642) );
  AOI22XL U4652 ( .A0(n6480), .A1(image_data[25]), .B0(n6479), .B1(
        image_data[153]), .Y(n5643) );
  AOI22XL U4653 ( .A0(n6450), .A1(image_data[97]), .B0(n6449), .B1(
        image_data[225]), .Y(n5628) );
  AOI22XL U4654 ( .A0(n6448), .A1(image_data[33]), .B0(n6447), .B1(
        image_data[161]), .Y(n5629) );
  AOI22XL U4655 ( .A0(n6446), .A1(image_data[65]), .B0(n6445), .B1(
        image_data[193]), .Y(n5630) );
  AOI22XL U4656 ( .A0(n6444), .A1(image_data[1]), .B0(n6443), .B1(
        image_data[129]), .Y(n5631) );
  AOI22XL U4657 ( .A0(n6458), .A1(image_data[81]), .B0(n6457), .B1(
        image_data[209]), .Y(n5634) );
  AOI22XL U4658 ( .A0(n6462), .A1(image_data[113]), .B0(n6461), .B1(
        image_data[241]), .Y(n5632) );
  AOI22XL U4659 ( .A0(n6460), .A1(image_data[49]), .B0(n6459), .B1(
        image_data[177]), .Y(n5633) );
  AOI22XL U4660 ( .A0(n6456), .A1(image_data[17]), .B0(n6455), .B1(
        image_data[145]), .Y(n5635) );
  NAND4XL U4661 ( .A(n5639), .B(n5638), .C(n5637), .D(n5636), .Y(n5645) );
  AOI22XL U4662 ( .A0(n6468), .A1(image_data[9]), .B0(n6467), .B1(
        image_data[137]), .Y(n5639) );
  AOI22XL U4663 ( .A0(n6470), .A1(image_data[73]), .B0(n6469), .B1(
        image_data[201]), .Y(n5638) );
  AOI22XL U4664 ( .A0(n6472), .A1(image_data[41]), .B0(n6471), .B1(
        image_data[169]), .Y(n5637) );
  AOI22XL U4665 ( .A0(n6550), .A1(image_data[111]), .B0(n6549), .B1(
        image_data[239]), .Y(n6551) );
  AOI22XL U4666 ( .A0(n6562), .A1(image_data[127]), .B0(n6561), .B1(
        image_data[255]), .Y(n6563) );
  AOI22XL U4667 ( .A0(n6538), .A1(image_data[119]), .B0(n6537), .B1(
        image_data[247]), .Y(n6539) );
  AOI22XL U4668 ( .A0(n6526), .A1(image_data[103]), .B0(n6525), .B1(
        image_data[231]), .Y(n6527) );
  AOI22XL U4669 ( .A0(n6550), .A1(image_data[367]), .B0(n6549), .B1(
        image_data[495]), .Y(n6507) );
  AOI22XL U4670 ( .A0(n6562), .A1(image_data[383]), .B0(n6561), .B1(
        image_data[511]), .Y(n6511) );
  AOI22XL U4671 ( .A0(n6538), .A1(image_data[375]), .B0(n6537), .B1(
        image_data[503]), .Y(n6503) );
  AOI22XL U4672 ( .A0(n6474), .A1(image_data[111]), .B0(n6473), .B1(
        image_data[239]), .Y(n6475) );
  AOI22XL U4673 ( .A0(n6462), .A1(image_data[119]), .B0(n6461), .B1(
        image_data[247]), .Y(n6463) );
  AOI22XL U4674 ( .A0(n6450), .A1(image_data[103]), .B0(n6449), .B1(
        image_data[231]), .Y(n6451) );
  AOI22XL U4675 ( .A0(n6486), .A1(image_data[127]), .B0(n6485), .B1(
        image_data[255]), .Y(n6487) );
  AOI22XL U4676 ( .A0(n6474), .A1(image_data[367]), .B0(n6473), .B1(
        image_data[495]), .Y(n6431) );
  AOI22XL U4677 ( .A0(n6462), .A1(image_data[375]), .B0(n6461), .B1(
        image_data[503]), .Y(n6427) );
  AOI22XL U4678 ( .A0(n6450), .A1(image_data[359]), .B0(n6449), .B1(
        image_data[487]), .Y(n6423) );
  AOI22XL U4679 ( .A0(n6474), .A1(image_data[364]), .B0(n6473), .B1(
        image_data[492]), .Y(n5718) );
  AOI22XL U4680 ( .A0(n6462), .A1(image_data[372]), .B0(n6461), .B1(
        image_data[500]), .Y(n5714) );
  AOI22XL U4681 ( .A0(n6450), .A1(image_data[356]), .B0(n6449), .B1(
        image_data[484]), .Y(n5710) );
  AOI22XL U4682 ( .A0(n6486), .A1(image_data[380]), .B0(n6485), .B1(
        image_data[508]), .Y(n5722) );
  AOI22XL U4683 ( .A0(n6538), .A1(image_data[116]), .B0(n6537), .B1(
        image_data[244]), .Y(n5776) );
  AOI22XL U4684 ( .A0(n6536), .A1(image_data[52]), .B0(n6535), .B1(
        image_data[180]), .Y(n5777) );
  AOI22XL U4685 ( .A0(n6534), .A1(image_data[84]), .B0(n6533), .B1(
        image_data[212]), .Y(n5778) );
  AOI22XL U4686 ( .A0(n6532), .A1(image_data[20]), .B0(n6531), .B1(
        image_data[148]), .Y(n5779) );
  AOI22XL U4687 ( .A0(n6526), .A1(image_data[100]), .B0(n6525), .B1(
        image_data[228]), .Y(n5772) );
  AOI22XL U4688 ( .A0(n6524), .A1(image_data[36]), .B0(n6523), .B1(
        image_data[164]), .Y(n5773) );
  AOI22XL U4689 ( .A0(n6522), .A1(image_data[68]), .B0(n6521), .B1(
        image_data[196]), .Y(n5774) );
  AOI22XL U4690 ( .A0(n6520), .A1(image_data[4]), .B0(n6519), .B1(
        image_data[132]), .Y(n5775) );
  AOI22XL U4691 ( .A0(n6562), .A1(image_data[124]), .B0(n6561), .B1(
        image_data[252]), .Y(n5784) );
  AOI22XL U4692 ( .A0(n6556), .A1(image_data[28]), .B0(n6555), .B1(
        image_data[156]), .Y(n5787) );
  AOI22XL U4693 ( .A0(n6560), .A1(image_data[60]), .B0(n6559), .B1(
        image_data[188]), .Y(n5785) );
  AOI22XL U4694 ( .A0(n6558), .A1(image_data[92]), .B0(n6557), .B1(
        image_data[220]), .Y(n5786) );
  NAND4XL U4695 ( .A(n5783), .B(n5782), .C(n5781), .D(n5780), .Y(n5789) );
  AOI22XL U4696 ( .A0(n6544), .A1(image_data[12]), .B0(n6543), .B1(
        image_data[140]), .Y(n5783) );
  AOI22XL U4697 ( .A0(n6546), .A1(image_data[76]), .B0(n6545), .B1(
        image_data[204]), .Y(n5782) );
  AOI22XL U4698 ( .A0(n6548), .A1(image_data[44]), .B0(n6547), .B1(
        image_data[172]), .Y(n5781) );
  AOI22XL U4699 ( .A0(n6538), .A1(image_data[372]), .B0(n6537), .B1(
        image_data[500]), .Y(n5756) );
  AOI22XL U4700 ( .A0(n6536), .A1(image_data[308]), .B0(n6535), .B1(
        image_data[436]), .Y(n5757) );
  AOI22XL U4701 ( .A0(n6534), .A1(image_data[340]), .B0(n6533), .B1(
        image_data[468]), .Y(n5758) );
  AOI22XL U4702 ( .A0(n6532), .A1(image_data[276]), .B0(n6531), .B1(
        image_data[404]), .Y(n5759) );
  AOI22XL U4703 ( .A0(n6526), .A1(image_data[356]), .B0(n6525), .B1(
        image_data[484]), .Y(n5752) );
  AOI22XL U4704 ( .A0(n6524), .A1(image_data[292]), .B0(n6523), .B1(
        image_data[420]), .Y(n5753) );
  AOI22XL U4705 ( .A0(n6522), .A1(image_data[324]), .B0(n6521), .B1(
        image_data[452]), .Y(n5754) );
  AOI22XL U4706 ( .A0(n6520), .A1(image_data[260]), .B0(n6519), .B1(
        image_data[388]), .Y(n5755) );
  AOI22XL U4707 ( .A0(n6562), .A1(image_data[380]), .B0(n6561), .B1(
        image_data[508]), .Y(n5764) );
  AOI22XL U4708 ( .A0(n6556), .A1(image_data[284]), .B0(n6555), .B1(
        image_data[412]), .Y(n5767) );
  AOI22XL U4709 ( .A0(n6560), .A1(image_data[316]), .B0(n6559), .B1(
        image_data[444]), .Y(n5765) );
  AOI22XL U4710 ( .A0(n6558), .A1(image_data[348]), .B0(n6557), .B1(
        image_data[476]), .Y(n5766) );
  NAND4XL U4711 ( .A(n5763), .B(n5762), .C(n5761), .D(n5760), .Y(n5769) );
  AOI22XL U4712 ( .A0(n6544), .A1(image_data[268]), .B0(n6543), .B1(
        image_data[396]), .Y(n5763) );
  AOI22XL U4713 ( .A0(n6546), .A1(image_data[332]), .B0(n6545), .B1(
        image_data[460]), .Y(n5762) );
  AOI22XL U4714 ( .A0(n6548), .A1(image_data[300]), .B0(n6547), .B1(
        image_data[428]), .Y(n5761) );
  AOI22XL U4715 ( .A0(n6462), .A1(image_data[116]), .B0(n6461), .B1(
        image_data[244]), .Y(n5734) );
  AOI22XL U4716 ( .A0(n6460), .A1(image_data[52]), .B0(n6459), .B1(
        image_data[180]), .Y(n5735) );
  AOI22XL U4717 ( .A0(n6458), .A1(image_data[84]), .B0(n6457), .B1(
        image_data[212]), .Y(n5736) );
  AOI22XL U4718 ( .A0(n6456), .A1(image_data[20]), .B0(n6455), .B1(
        image_data[148]), .Y(n5737) );
  AOI22XL U4719 ( .A0(n6450), .A1(image_data[100]), .B0(n6449), .B1(
        image_data[228]), .Y(n5730) );
  AOI22XL U4720 ( .A0(n6448), .A1(image_data[36]), .B0(n6447), .B1(
        image_data[164]), .Y(n5731) );
  AOI22XL U4721 ( .A0(n6446), .A1(image_data[68]), .B0(n6445), .B1(
        image_data[196]), .Y(n5732) );
  AOI22XL U4722 ( .A0(n6444), .A1(image_data[4]), .B0(n6443), .B1(
        image_data[132]), .Y(n5733) );
  AOI22XL U4723 ( .A0(n6486), .A1(image_data[124]), .B0(n6485), .B1(
        image_data[252]), .Y(n5742) );
  AOI22XL U4724 ( .A0(n6484), .A1(image_data[60]), .B0(n6483), .B1(
        image_data[188]), .Y(n5743) );
  AOI22XL U4725 ( .A0(n6482), .A1(image_data[92]), .B0(n6481), .B1(
        image_data[220]), .Y(n5744) );
  AOI22XL U4726 ( .A0(n6480), .A1(image_data[28]), .B0(n6479), .B1(
        image_data[156]), .Y(n5745) );
  NAND4XL U4727 ( .A(n5741), .B(n5740), .C(n5739), .D(n5738), .Y(n5747) );
  AOI22XL U4728 ( .A0(n6468), .A1(image_data[12]), .B0(n6467), .B1(
        image_data[140]), .Y(n5741) );
  AOI22XL U4729 ( .A0(n6470), .A1(image_data[76]), .B0(n6469), .B1(
        image_data[204]), .Y(n5740) );
  AOI22XL U4730 ( .A0(n6472), .A1(image_data[44]), .B0(n6471), .B1(
        image_data[172]), .Y(n5739) );
  AOI22XL U4731 ( .A0(n6474), .A1(image_data[106]), .B0(n6473), .B1(
        image_data[234]), .Y(n5069) );
  AOI22XL U4732 ( .A0(n6474), .A1(image_data[362]), .B0(n6473), .B1(
        image_data[490]), .Y(n5038) );
  OAI211X1 U4733 ( .A0(n4977), .A1(n5120), .B0(n4976), .C0(n4975), .Y(n5007)
         );
  AOI22XL U4734 ( .A0(n5117), .A1(n4876), .B0(N2780), .B1(n5115), .Y(n4977) );
  AOI22XL U4735 ( .A0(n5096), .A1(n4974), .B0(n5124), .B1(n4973), .Y(n4975) );
  AOI22XL U4736 ( .A0(n5149), .A1(n4996), .B0(n5148), .B1(n4995), .Y(n4999) );
  AOI21XL U4737 ( .A0(n5131), .A1(n4982), .B0(n5129), .Y(n4983) );
  AOI22XL U4738 ( .A0(n6550), .A1(image_data[106]), .B0(n6549), .B1(
        image_data[234]), .Y(n5241) );
  AOI22XL U4739 ( .A0(n6562), .A1(image_data[122]), .B0(n6561), .B1(
        image_data[250]), .Y(n5245) );
  AOI22XL U4740 ( .A0(n6526), .A1(image_data[98]), .B0(n6525), .B1(
        image_data[226]), .Y(n5233) );
  AOI22XL U4741 ( .A0(n6534), .A1(image_data[82]), .B0(n6533), .B1(
        image_data[210]), .Y(n5239) );
  AOI22XL U4742 ( .A0(n6550), .A1(image_data[362]), .B0(n6549), .B1(
        image_data[490]), .Y(n5210) );
  AOI22XL U4743 ( .A0(n6562), .A1(image_data[378]), .B0(n6561), .B1(
        image_data[506]), .Y(n5225) );
  AOI22XL U4744 ( .A0(n6526), .A1(image_data[354]), .B0(n6525), .B1(
        image_data[482]), .Y(n5198) );
  AOI22XL U4745 ( .A0(n3935), .A1(image_data[370]), .B0(n3888), .B1(
        image_data[498]), .Y(n3775) );
  AOI22XL U4746 ( .A0(n3887), .A1(image_data[306]), .B0(n3936), .B1(
        image_data[434]), .Y(n3776) );
  AOI22XL U4747 ( .A0(n3884), .A1(image_data[274]), .B0(n3934), .B1(
        image_data[402]), .Y(n3778) );
  AOI22XL U4748 ( .A0(n3885), .A1(image_data[338]), .B0(n3886), .B1(
        image_data[466]), .Y(n3777) );
  NAND4XL U4749 ( .A(n3796), .B(n3795), .C(n3794), .D(n3793), .Y(n3819) );
  AOI22XL U4750 ( .A0(n3791), .A1(image_data[34]), .B0(n3929), .B1(
        image_data[162]), .Y(n3794) );
  AOI22XL U4751 ( .A0(n3897), .A1(image_data[2]), .B0(n3896), .B1(
        image_data[130]), .Y(n3796) );
  AOI22XL U4752 ( .A0(n3893), .A1(image_data[98]), .B0(n3792), .B1(
        image_data[226]), .Y(n3793) );
  NAND4XL U4753 ( .A(n3815), .B(n3814), .C(n3813), .D(n3812), .Y(n3816) );
  AOI22XL U4754 ( .A0(n3875), .A1(image_data[90]), .B0(n3810), .B1(
        image_data[218]), .Y(n3814) );
  AOI22XL U4755 ( .A0(n3877), .A1(image_data[58]), .B0(n3949), .B1(
        image_data[186]), .Y(n3813) );
  AOI22XL U4756 ( .A0(n3874), .A1(image_data[26]), .B0(n3948), .B1(
        image_data[154]), .Y(n3815) );
  NAND4XL U4757 ( .A(n3809), .B(n3808), .C(n3807), .D(n3806), .Y(n3817) );
  AOI22XL U4758 ( .A0(n3866), .A1(image_data[74]), .B0(n3804), .B1(
        image_data[202]), .Y(n3808) );
  AOI22XL U4759 ( .A0(n3865), .A1(image_data[10]), .B0(n3941), .B1(
        image_data[138]), .Y(n3809) );
  AOI22XL U4760 ( .A0(n3942), .A1(image_data[42]), .B0(n3943), .B1(
        image_data[170]), .Y(n3807) );
  NAND4XL U4761 ( .A(n3803), .B(n3802), .C(n3801), .D(n3800), .Y(n3818) );
  AOI22XL U4762 ( .A0(n3885), .A1(image_data[82]), .B0(n3797), .B1(
        image_data[210]), .Y(n3802) );
  AOI22XL U4763 ( .A0(n3884), .A1(image_data[18]), .B0(n3934), .B1(
        image_data[146]), .Y(n3803) );
  AOI22XL U4764 ( .A0(n3798), .A1(image_data[50]), .B0(n3936), .B1(
        image_data[178]), .Y(n3801) );
  NAND4XL U4765 ( .A(n3774), .B(n3773), .C(n3772), .D(n3771), .Y(n3790) );
  AOI22XL U4766 ( .A0(n3928), .A1(image_data[290]), .B0(n3929), .B1(
        image_data[418]), .Y(n3772) );
  AOI22XL U4767 ( .A0(n3897), .A1(image_data[258]), .B0(n3896), .B1(
        image_data[386]), .Y(n3774) );
  AOI22XL U4768 ( .A0(n3893), .A1(image_data[354]), .B0(n3894), .B1(
        image_data[482]), .Y(n3771) );
  NAND4XL U4769 ( .A(n3786), .B(n3785), .C(n3784), .D(n3783), .Y(n3787) );
  AOI22XL U4770 ( .A0(n3875), .A1(image_data[346]), .B0(n3876), .B1(
        image_data[474]), .Y(n3785) );
  AOI22XL U4771 ( .A0(n3877), .A1(image_data[314]), .B0(n3949), .B1(
        image_data[442]), .Y(n3784) );
  AOI22XL U4772 ( .A0(n3874), .A1(image_data[282]), .B0(n3948), .B1(
        image_data[410]), .Y(n3786) );
  NAND4XL U4773 ( .A(n3782), .B(n3781), .C(n3780), .D(n3779), .Y(n3788) );
  AOI22XL U4774 ( .A0(n3866), .A1(image_data[330]), .B0(n3867), .B1(
        image_data[458]), .Y(n3781) );
  AOI22XL U4775 ( .A0(n3865), .A1(image_data[266]), .B0(n3941), .B1(
        image_data[394]), .Y(n3782) );
  AOI22XL U4776 ( .A0(n3942), .A1(image_data[298]), .B0(n3943), .B1(
        image_data[426]), .Y(n3780) );
  AOI22XL U4777 ( .A0(n3895), .A1(image_data[122]), .B0(n3364), .B1(
        image_data[250]), .Y(n3854) );
  AOI22XL U4778 ( .A0(n3888), .A1(image_data[42]), .B0(n3935), .B1(
        image_data[170]), .Y(n3851) );
  AOI22XL U4779 ( .A0(n3869), .A1(image_data[34]), .B0(n3868), .B1(
        image_data[162]), .Y(n3843) );
  AOI22XL U4780 ( .A0(n3879), .A1(image_data[50]), .B0(n3878), .B1(
        image_data[178]), .Y(n3847) );
  AOI22XL U4781 ( .A0(n3895), .A1(image_data[378]), .B0(n3364), .B1(
        image_data[506]), .Y(n3834) );
  AOI22XL U4782 ( .A0(n3888), .A1(image_data[298]), .B0(n3935), .B1(
        image_data[426]), .Y(n3831) );
  AOI22XL U4783 ( .A0(n3869), .A1(image_data[290]), .B0(n3868), .B1(
        image_data[418]), .Y(n3823) );
  AOI22XL U4784 ( .A0(n3895), .A1(image_data[69]), .B0(n3364), .B1(
        image_data[197]), .Y(n4515) );
  AOI22XL U4785 ( .A0(n3878), .A1(image_data[125]), .B0(n3879), .B1(
        image_data[253]), .Y(n4525) );
  AOI22XL U4786 ( .A0(n3868), .A1(image_data[109]), .B0(n3869), .B1(
        image_data[237]), .Y(n4521) );
  AOI22XL U4787 ( .A0(n3935), .A1(image_data[117]), .B0(n3888), .B1(
        image_data[245]), .Y(n4517) );
  AOI22XL U4788 ( .A0(n3895), .A1(image_data[325]), .B0(n3364), .B1(
        image_data[453]), .Y(n4495) );
  AOI22XL U4789 ( .A0(n3878), .A1(image_data[381]), .B0(n3879), .B1(
        image_data[509]), .Y(n4505) );
  AOI22XL U4790 ( .A0(n3868), .A1(image_data[365]), .B0(n3869), .B1(
        image_data[493]), .Y(n4501) );
  AOI22XL U4791 ( .A0(n3895), .A1(image_data[125]), .B0(n3364), .B1(
        image_data[253]), .Y(n3550) );
  AOI22XL U4792 ( .A0(n3888), .A1(image_data[45]), .B0(n3935), .B1(
        image_data[173]), .Y(n3547) );
  AOI22XL U4793 ( .A0(n3879), .A1(image_data[53]), .B0(n3878), .B1(
        image_data[181]), .Y(n3543) );
  AOI22XL U4794 ( .A0(n3869), .A1(image_data[37]), .B0(n3868), .B1(
        image_data[165]), .Y(n3539) );
  AOI22XL U4795 ( .A0(n3895), .A1(image_data[381]), .B0(n3364), .B1(
        image_data[509]), .Y(n3530) );
  AOI22XL U4796 ( .A0(n3888), .A1(image_data[301]), .B0(n3935), .B1(
        image_data[429]), .Y(n3527) );
  AOI22XL U4797 ( .A0(n3879), .A1(image_data[309]), .B0(n3878), .B1(
        image_data[437]), .Y(n3523) );
  AOI22XL U4798 ( .A0(n3878), .A1(image_data[124]), .B0(n3879), .B1(
        image_data[252]), .Y(n4483) );
  AOI22XL U4799 ( .A0(n3868), .A1(image_data[108]), .B0(n3869), .B1(
        image_data[236]), .Y(n4479) );
  AOI22XL U4800 ( .A0(n3893), .A1(image_data[100]), .B0(n3894), .B1(
        image_data[228]), .Y(n4471) );
  AOI22XL U4801 ( .A0(n3935), .A1(image_data[116]), .B0(n3888), .B1(
        image_data[244]), .Y(n4475) );
  AOI22XL U4802 ( .A0(n3878), .A1(image_data[380]), .B0(n3879), .B1(
        image_data[508]), .Y(n4463) );
  AOI22XL U4803 ( .A0(n3868), .A1(image_data[364]), .B0(n3869), .B1(
        image_data[492]), .Y(n4459) );
  AOI22XL U4804 ( .A0(n3893), .A1(image_data[356]), .B0(n3894), .B1(
        image_data[484]), .Y(n4451) );
  AOI22XL U4805 ( .A0(n3895), .A1(image_data[124]), .B0(n3364), .B1(
        image_data[252]), .Y(n3676) );
  AOI22XL U4806 ( .A0(n3888), .A1(image_data[44]), .B0(n3935), .B1(
        image_data[172]), .Y(n3673) );
  AOI22XL U4807 ( .A0(n3869), .A1(image_data[36]), .B0(n3868), .B1(
        image_data[164]), .Y(n3665) );
  AOI22XL U4808 ( .A0(n3879), .A1(image_data[52]), .B0(n3878), .B1(
        image_data[180]), .Y(n3669) );
  AOI22XL U4809 ( .A0(n3888), .A1(image_data[300]), .B0(n3935), .B1(
        image_data[428]), .Y(n3653) );
  AOI22XL U4810 ( .A0(n3869), .A1(image_data[292]), .B0(n3868), .B1(
        image_data[420]), .Y(n3645) );
  AOI22XL U4811 ( .A0(n3879), .A1(image_data[308]), .B0(n3878), .B1(
        image_data[436]), .Y(n3649) );
  AOI22XL U4812 ( .A0(n6550), .A1(image_data[109]), .B0(n6549), .B1(
        image_data[237]), .Y(n6001) );
  AOI22XL U4813 ( .A0(n6538), .A1(image_data[117]), .B0(n6537), .B1(
        image_data[245]), .Y(n5997) );
  AOI22XL U4814 ( .A0(n6526), .A1(image_data[101]), .B0(n6525), .B1(
        image_data[229]), .Y(n5993) );
  AOI22XL U4815 ( .A0(n6562), .A1(image_data[125]), .B0(n6561), .B1(
        image_data[253]), .Y(n6005) );
  AOI22XL U4816 ( .A0(n6550), .A1(image_data[365]), .B0(n6549), .B1(
        image_data[493]), .Y(n5981) );
  AOI22XL U4817 ( .A0(n6538), .A1(image_data[373]), .B0(n6537), .B1(
        image_data[501]), .Y(n5977) );
  AOI22XL U4818 ( .A0(n6526), .A1(image_data[357]), .B0(n6525), .B1(
        image_data[485]), .Y(n5973) );
  AOI22XL U4819 ( .A0(n6474), .A1(image_data[109]), .B0(n6473), .B1(
        image_data[237]), .Y(n5959) );
  AOI22XL U4820 ( .A0(n6462), .A1(image_data[117]), .B0(n6461), .B1(
        image_data[245]), .Y(n5955) );
  AOI22XL U4821 ( .A0(n6450), .A1(image_data[101]), .B0(n6449), .B1(
        image_data[229]), .Y(n5951) );
  AOI22XL U4822 ( .A0(n6486), .A1(image_data[125]), .B0(n6485), .B1(
        image_data[253]), .Y(n5963) );
  AOI22XL U4823 ( .A0(n6474), .A1(image_data[365]), .B0(n6473), .B1(
        image_data[493]), .Y(n5939) );
  AOI22XL U4824 ( .A0(n6462), .A1(image_data[373]), .B0(n6461), .B1(
        image_data[501]), .Y(n5935) );
  AOI22XL U4825 ( .A0(n6450), .A1(image_data[357]), .B0(n6449), .B1(
        image_data[485]), .Y(n5931) );
  AOI22XL U4826 ( .A0(n3895), .A1(image_data[70]), .B0(n3364), .B1(
        image_data[198]), .Y(n4425) );
  AOI22XL U4827 ( .A0(n3878), .A1(image_data[126]), .B0(n3879), .B1(
        image_data[254]), .Y(n4441) );
  AOI22XL U4828 ( .A0(n3868), .A1(image_data[110]), .B0(n3869), .B1(
        image_data[238]), .Y(n4435) );
  NOR2XL U4829 ( .A(n3484), .B(n3471), .Y(n4427) );
  NOR2XL U4830 ( .A(n3487), .B(n3471), .Y(n4428) );
  AOI22XL U4831 ( .A0(n3935), .A1(image_data[118]), .B0(n3888), .B1(
        image_data[246]), .Y(n4429) );
  NOR2XL U4832 ( .A(n5002), .B(n3487), .Y(n4422) );
  AOI22XL U4833 ( .A0(n3895), .A1(image_data[326]), .B0(n3364), .B1(
        image_data[454]), .Y(n4404) );
  NOR2XL U4834 ( .A(n3487), .B(n4588), .Y(n4440) );
  NOR2XL U4835 ( .A(n3484), .B(n4588), .Y(n4439) );
  AOI22XL U4836 ( .A0(n3878), .A1(image_data[382]), .B0(n3879), .B1(
        image_data[510]), .Y(n4414) );
  NOR2XL U4837 ( .A(n3487), .B(n3476), .Y(n4434) );
  AOI22XL U4838 ( .A0(n3868), .A1(image_data[366]), .B0(n3869), .B1(
        image_data[494]), .Y(n4410) );
  AOI22XL U4839 ( .A0(n3895), .A1(image_data[126]), .B0(n3364), .B1(
        image_data[254]), .Y(n4055) );
  AOI22XL U4840 ( .A0(n3888), .A1(image_data[46]), .B0(n3935), .B1(
        image_data[174]), .Y(n4052) );
  AOI22XL U4841 ( .A0(n3879), .A1(image_data[54]), .B0(n3878), .B1(
        image_data[182]), .Y(n4048) );
  AOI22XL U4842 ( .A0(n3869), .A1(image_data[38]), .B0(n3868), .B1(
        image_data[166]), .Y(n4044) );
  AOI22XL U4843 ( .A0(n3895), .A1(image_data[382]), .B0(n3364), .B1(
        image_data[510]), .Y(n4035) );
  AOI22XL U4844 ( .A0(n3888), .A1(image_data[302]), .B0(n3935), .B1(
        image_data[430]), .Y(n4032) );
  AOI22XL U4845 ( .A0(n3879), .A1(image_data[310]), .B0(n3878), .B1(
        image_data[438]), .Y(n4028) );
  AOI22XL U4846 ( .A0(n3895), .A1(image_data[59]), .B0(n3364), .B1(
        image_data[187]), .Y(n4309) );
  AOI22XL U4847 ( .A0(n3935), .A1(image_data[107]), .B0(n3888), .B1(
        image_data[235]), .Y(n4304) );
  AOI22XL U4848 ( .A0(n4721), .A1(image_data[115]), .B0(n3879), .B1(
        image_data[243]), .Y(n4300) );
  AOI22XL U4849 ( .A0(n4714), .A1(image_data[99]), .B0(n3869), .B1(
        image_data[227]), .Y(n4296) );
  AOI22XL U4850 ( .A0(n3895), .A1(image_data[315]), .B0(n3364), .B1(
        image_data[443]), .Y(n4289) );
  AOI22XL U4851 ( .A0(n3868), .A1(image_data[355]), .B0(n3869), .B1(
        image_data[483]), .Y(n4276) );
  AOI22XL U4852 ( .A0(n3935), .A1(image_data[363]), .B0(n3888), .B1(
        image_data[491]), .Y(n4284) );
  AOI22XL U4853 ( .A0(n3364), .A1(image_data[3]), .B0(n3895), .B1(
        image_data[131]), .Y(n4088) );
  AOI22XL U4854 ( .A0(n3874), .A1(image_data[91]), .B0(n3948), .B1(
        image_data[219]), .Y(n4099) );
  AOI22XL U4855 ( .A0(n3869), .A1(image_data[43]), .B0(n3868), .B1(
        image_data[171]), .Y(n4094) );
  AOI22XL U4856 ( .A0(n3884), .A1(image_data[83]), .B0(n3934), .B1(
        image_data[211]), .Y(n4091) );
  AOI22XL U4857 ( .A0(n3364), .A1(image_data[259]), .B0(n3895), .B1(
        image_data[387]), .Y(n4068) );
  AOI22XL U4858 ( .A0(n3874), .A1(image_data[347]), .B0(n3948), .B1(
        image_data[475]), .Y(n4079) );
  AOI22XL U4859 ( .A0(n3942), .A1(image_data[363]), .B0(n3943), .B1(
        image_data[491]), .Y(n4073) );
  AOI22XL U4860 ( .A0(n3884), .A1(image_data[339]), .B0(n3934), .B1(
        image_data[467]), .Y(n4071) );
  AOI22XL U4861 ( .A0(n3895), .A1(image_data[60]), .B0(n3364), .B1(
        image_data[188]), .Y(n4267) );
  AOI22XL U4862 ( .A0(n3878), .A1(image_data[116]), .B0(n3879), .B1(
        image_data[244]), .Y(n4258) );
  AOI22XL U4863 ( .A0(n3868), .A1(image_data[100]), .B0(n3869), .B1(
        image_data[228]), .Y(n4254) );
  AOI22XL U4864 ( .A0(n3935), .A1(image_data[108]), .B0(n3888), .B1(
        image_data[236]), .Y(n4262) );
  AOI22XL U4865 ( .A0(n3895), .A1(image_data[316]), .B0(n3364), .B1(
        image_data[444]), .Y(n4247) );
  AOI22XL U4866 ( .A0(n3878), .A1(image_data[372]), .B0(n3879), .B1(
        image_data[500]), .Y(n4238) );
  AOI22XL U4867 ( .A0(n3868), .A1(image_data[356]), .B0(n3869), .B1(
        image_data[484]), .Y(n4234) );
  AOI22XL U4868 ( .A0(n3879), .A1(image_data[60]), .B0(n3878), .B1(
        image_data[188]), .Y(n4183) );
  AOI22XL U4869 ( .A0(n3869), .A1(image_data[44]), .B0(n3868), .B1(
        image_data[172]), .Y(n4179) );
  AOI22XL U4870 ( .A0(n3894), .A1(image_data[36]), .B0(n3893), .B1(
        image_data[164]), .Y(n4171) );
  AOI22XL U4871 ( .A0(n3888), .A1(image_data[52]), .B0(n3935), .B1(
        image_data[180]), .Y(n4175) );
  AOI22XL U4872 ( .A0(n3879), .A1(image_data[316]), .B0(n3878), .B1(
        image_data[444]), .Y(n4163) );
  AOI22XL U4873 ( .A0(n3869), .A1(image_data[300]), .B0(n3868), .B1(
        image_data[428]), .Y(n4159) );
  AOI22XL U4874 ( .A0(n3894), .A1(image_data[292]), .B0(n3893), .B1(
        image_data[420]), .Y(n4151) );
  AOI22XL U4875 ( .A0(n3895), .A1(image_data[56]), .B0(n3364), .B1(
        image_data[184]), .Y(n4819) );
  AOI22XL U4876 ( .A0(n3935), .A1(image_data[104]), .B0(n3888), .B1(
        image_data[232]), .Y(n4814) );
  AOI22XL U4877 ( .A0(n3874), .A1(image_data[16]), .B0(n3948), .B1(
        image_data[144]), .Y(n4813) );
  AOI22XL U4878 ( .A0(n3942), .A1(image_data[32]), .B0(n3943), .B1(
        image_data[160]), .Y(n4807) );
  AOI22XL U4879 ( .A0(n3895), .A1(image_data[312]), .B0(n3364), .B1(
        image_data[440]), .Y(n4799) );
  AOI22XL U4880 ( .A0(n3935), .A1(image_data[360]), .B0(n3888), .B1(
        image_data[488]), .Y(n4794) );
  AOI22XL U4881 ( .A0(n3874), .A1(image_data[272]), .B0(n3948), .B1(
        image_data[400]), .Y(n4793) );
  AOI22XL U4882 ( .A0(n3874), .A1(image_data[344]), .B0(n3948), .B1(
        image_data[472]), .Y(n4610) );
  AOI22XL U4883 ( .A0(n3942), .A1(image_data[360]), .B0(n3943), .B1(
        image_data[488]), .Y(n4604) );
  AOI22XL U4884 ( .A0(n3884), .A1(image_data[336]), .B0(n3934), .B1(
        image_data[464]), .Y(n4602) );
  AOI22XL U4885 ( .A0(n3928), .A1(image_data[352]), .B0(n3929), .B1(
        image_data[480]), .Y(n4596) );
  AOI22XL U4886 ( .A0(n3874), .A1(image_data[88]), .B0(n3948), .B1(
        image_data[216]), .Y(n4630) );
  AOI22XL U4887 ( .A0(n3877), .A1(image_data[120]), .B0(n3949), .B1(
        image_data[248]), .Y(n4628) );
  AOI22XL U4888 ( .A0(n3879), .A1(image_data[56]), .B0(n4721), .B1(
        image_data[184]), .Y(n4629) );
  AOI22XL U4889 ( .A0(n3876), .A1(image_data[24]), .B0(n4719), .B1(
        image_data[152]), .Y(n4631) );
  AOI22XL U4890 ( .A0(n3942), .A1(image_data[104]), .B0(n3943), .B1(
        image_data[232]), .Y(n4624) );
  AOI22XL U4891 ( .A0(n3865), .A1(image_data[72]), .B0(n3941), .B1(
        image_data[200]), .Y(n4626) );
  AOI22XL U4892 ( .A0(n3869), .A1(image_data[40]), .B0(n4714), .B1(
        image_data[168]), .Y(n4625) );
  AOI22XL U4893 ( .A0(n3867), .A1(image_data[8]), .B0(n4713), .B1(
        image_data[136]), .Y(n4627) );
  AOI22XL U4894 ( .A0(n3884), .A1(image_data[80]), .B0(n3934), .B1(
        image_data[208]), .Y(n4622) );
  AOI22XL U4895 ( .A0(n3888), .A1(image_data[48]), .B0(n3935), .B1(
        image_data[176]), .Y(n4621) );
  AOI22XL U4896 ( .A0(n3887), .A1(image_data[112]), .B0(n3936), .B1(
        image_data[240]), .Y(n4620) );
  AOI22XL U4897 ( .A0(n3886), .A1(image_data[16]), .B0(n4707), .B1(
        image_data[144]), .Y(n4623) );
  NAND4XL U4898 ( .A(n4619), .B(n4618), .C(n4617), .D(n4616), .Y(n4635) );
  AOI22XL U4899 ( .A0(n3897), .A1(image_data[64]), .B0(n3896), .B1(
        image_data[192]), .Y(n4618) );
  AOI22XL U4900 ( .A0(n3928), .A1(image_data[96]), .B0(n3929), .B1(
        image_data[224]), .Y(n4616) );
  AOI22XL U4901 ( .A0(n3894), .A1(image_data[32]), .B0(n3893), .B1(
        image_data[160]), .Y(n4617) );
  AOI22XL U4902 ( .A0(n3895), .A1(image_data[123]), .B0(n3364), .B1(
        image_data[251]), .Y(n4140) );
  AOI22XL U4903 ( .A0(n3888), .A1(image_data[43]), .B0(n3935), .B1(
        image_data[171]), .Y(n4137) );
  AOI22XL U4904 ( .A0(n3869), .A1(image_data[35]), .B0(n3868), .B1(
        image_data[163]), .Y(n4129) );
  AOI22XL U4905 ( .A0(n3879), .A1(image_data[51]), .B0(n3878), .B1(
        image_data[179]), .Y(n4133) );
  AOI22XL U4906 ( .A0(n3895), .A1(image_data[379]), .B0(n3364), .B1(
        image_data[507]), .Y(n4120) );
  AOI22XL U4907 ( .A0(n3888), .A1(image_data[299]), .B0(n3935), .B1(
        image_data[427]), .Y(n4117) );
  AOI22XL U4908 ( .A0(n3869), .A1(image_data[291]), .B0(n3868), .B1(
        image_data[419]), .Y(n4109) );
  AOI22XL U4909 ( .A0(n3895), .A1(image_data[61]), .B0(n3364), .B1(
        image_data[189]), .Y(n4225) );
  AOI22XL U4910 ( .A0(n3935), .A1(image_data[109]), .B0(n3888), .B1(
        image_data[237]), .Y(n4220) );
  AOI22XL U4911 ( .A0(n4720), .A1(image_data[21]), .B0(n3948), .B1(
        image_data[149]), .Y(n4219) );
  AOI22XL U4912 ( .A0(n3942), .A1(image_data[37]), .B0(n3943), .B1(
        image_data[165]), .Y(n4213) );
  AOI22XL U4913 ( .A0(n3895), .A1(image_data[317]), .B0(n3364), .B1(
        image_data[445]), .Y(n4205) );
  AOI22XL U4914 ( .A0(n3878), .A1(image_data[373]), .B0(n3879), .B1(
        image_data[501]), .Y(n4196) );
  AOI22XL U4915 ( .A0(n3868), .A1(image_data[357]), .B0(n3869), .B1(
        image_data[485]), .Y(n4192) );
  AOI22XL U4916 ( .A0(n3879), .A1(image_data[61]), .B0(n3878), .B1(
        image_data[189]), .Y(n4014) );
  AOI22XL U4917 ( .A0(n3869), .A1(image_data[45]), .B0(n3868), .B1(
        image_data[173]), .Y(n4010) );
  AOI22XL U4918 ( .A0(n3894), .A1(image_data[37]), .B0(n3893), .B1(
        image_data[165]), .Y(n4002) );
  AOI22XL U4919 ( .A0(n3884), .A1(image_data[85]), .B0(n3934), .B1(
        image_data[213]), .Y(n4007) );
  AOI22XL U4920 ( .A0(n3879), .A1(image_data[317]), .B0(n3878), .B1(
        image_data[445]), .Y(n3994) );
  AOI22XL U4921 ( .A0(n3869), .A1(image_data[301]), .B0(n3868), .B1(
        image_data[429]), .Y(n3990) );
  AOI22XL U4922 ( .A0(n3364), .A1(image_data[261]), .B0(n3895), .B1(
        image_data[389]), .Y(n3984) );
  AOI22XL U4923 ( .A0(n3895), .A1(image_data[62]), .B0(n3364), .B1(
        image_data[190]), .Y(n4351) );
  AOI22XL U4924 ( .A0(n3884), .A1(image_data[14]), .B0(n3934), .B1(
        image_data[142]), .Y(n4349) );
  AOI22XL U4925 ( .A0(n3874), .A1(image_data[22]), .B0(n3948), .B1(
        image_data[150]), .Y(n4345) );
  AOI22XL U4926 ( .A0(n3942), .A1(image_data[38]), .B0(n3943), .B1(
        image_data[166]), .Y(n4339) );
  AOI22XL U4927 ( .A0(n3895), .A1(image_data[318]), .B0(n3364), .B1(
        image_data[446]), .Y(n4331) );
  AOI22XL U4928 ( .A0(n3884), .A1(image_data[270]), .B0(n3934), .B1(
        image_data[398]), .Y(n4329) );
  AOI22XL U4929 ( .A0(n3874), .A1(image_data[278]), .B0(n3948), .B1(
        image_data[406]), .Y(n4325) );
  AOI22XL U4930 ( .A0(n3874), .A1(image_data[94]), .B0(n3948), .B1(
        image_data[222]), .Y(n3720) );
  AOI22XL U4931 ( .A0(n4754), .A1(image_data[110]), .B0(n3943), .B1(
        image_data[238]), .Y(n3714) );
  AOI22XL U4932 ( .A0(n3894), .A1(image_data[38]), .B0(n3893), .B1(
        image_data[166]), .Y(n3707) );
  AOI22XL U4933 ( .A0(n3884), .A1(image_data[86]), .B0(n3934), .B1(
        image_data[214]), .Y(n3712) );
  AOI22XL U4934 ( .A0(n3874), .A1(image_data[350]), .B0(n3948), .B1(
        image_data[478]), .Y(n3700) );
  AOI22XL U4935 ( .A0(n4754), .A1(image_data[366]), .B0(n3943), .B1(
        image_data[494]), .Y(n3694) );
  AOI22XL U4936 ( .A0(n3894), .A1(image_data[294]), .B0(n3893), .B1(
        image_data[422]), .Y(n3687) );
  AOI22XL U4937 ( .A0(n3884), .A1(image_data[342]), .B0(n3934), .B1(
        image_data[470]), .Y(n3692) );
  AOI22XL U4938 ( .A0(n3878), .A1(image_data[127]), .B0(n3879), .B1(
        image_data[255]), .Y(n3592) );
  AOI22XL U4939 ( .A0(n3868), .A1(image_data[111]), .B0(n3869), .B1(
        image_data[239]), .Y(n3588) );
  AOI22XL U4940 ( .A0(n3893), .A1(image_data[103]), .B0(n3894), .B1(
        image_data[231]), .Y(n3580) );
  AOI22XL U4941 ( .A0(n3935), .A1(image_data[119]), .B0(n3888), .B1(
        image_data[247]), .Y(n3584) );
  AOI22XL U4942 ( .A0(n3878), .A1(image_data[383]), .B0(n3879), .B1(
        image_data[511]), .Y(n3572) );
  NOR2X1 U4943 ( .A(n3484), .B(n3476), .Y(n4433) );
  AOI22XL U4944 ( .A0(n3868), .A1(image_data[367]), .B0(n3869), .B1(
        image_data[495]), .Y(n3568) );
  AOI22XL U4945 ( .A0(n3893), .A1(image_data[359]), .B0(n3894), .B1(
        image_data[487]), .Y(n3560) );
  AOI22XL U4946 ( .A0(n3895), .A1(image_data[127]), .B0(n3364), .B1(
        image_data[255]), .Y(n3634) );
  AOI22XL U4947 ( .A0(n3888), .A1(image_data[47]), .B0(n3935), .B1(
        image_data[175]), .Y(n3631) );
  AOI22XL U4948 ( .A0(n3879), .A1(image_data[55]), .B0(n3878), .B1(
        image_data[183]), .Y(n3627) );
  AOI22XL U4949 ( .A0(n3869), .A1(image_data[39]), .B0(n3868), .B1(
        image_data[167]), .Y(n3623) );
  AOI22XL U4950 ( .A0(n3894), .A1(image_data[287]), .B0(n3893), .B1(
        image_data[415]), .Y(n3617) );
  AOI22XL U4951 ( .A0(n3888), .A1(image_data[303]), .B0(n3935), .B1(
        image_data[431]), .Y(n3611) );
  AOI22XL U4952 ( .A0(n3879), .A1(image_data[311]), .B0(n3878), .B1(
        image_data[439]), .Y(n3607) );
  AOI22XL U4953 ( .A0(n3895), .A1(image_data[58]), .B0(n3364), .B1(
        image_data[186]), .Y(n3919) );
  AOI22XL U4954 ( .A0(n3887), .A1(image_data[42]), .B0(n3936), .B1(
        image_data[170]), .Y(n3915) );
  AOI22XL U4955 ( .A0(n3878), .A1(image_data[114]), .B0(n3879), .B1(
        image_data[242]), .Y(n3910) );
  AOI22XL U4956 ( .A0(n3942), .A1(image_data[34]), .B0(n3943), .B1(
        image_data[162]), .Y(n3907) );
  AOI22XL U4957 ( .A0(n3895), .A1(image_data[314]), .B0(n3364), .B1(
        image_data[442]), .Y(n3899) );
  AOI22XL U4958 ( .A0(n3887), .A1(image_data[298]), .B0(n3936), .B1(
        image_data[426]), .Y(n3890) );
  AOI22XL U4959 ( .A0(n3874), .A1(image_data[274]), .B0(n3948), .B1(
        image_data[402]), .Y(n3883) );
  AOI22XL U4960 ( .A0(n3364), .A1(image_data[2]), .B0(n3895), .B1(
        image_data[130]), .Y(n3961) );
  AOI22XL U4961 ( .A0(n3874), .A1(image_data[90]), .B0(n3948), .B1(
        image_data[218]), .Y(n3972) );
  AOI22XL U4962 ( .A0(n3942), .A1(image_data[106]), .B0(n3943), .B1(
        image_data[234]), .Y(n3966) );
  AOI22XL U4963 ( .A0(n3884), .A1(image_data[82]), .B0(n3934), .B1(
        image_data[210]), .Y(n3964) );
  AOI22XL U4964 ( .A0(n3874), .A1(image_data[346]), .B0(n3948), .B1(
        image_data[474]), .Y(n3952) );
  AOI22XL U4965 ( .A0(n3942), .A1(image_data[362]), .B0(n3943), .B1(
        image_data[490]), .Y(n3944) );
  AOI22XL U4966 ( .A0(n3884), .A1(image_data[338]), .B0(n3934), .B1(
        image_data[466]), .Y(n3939) );
  AOI22XL U4967 ( .A0(n3928), .A1(image_data[354]), .B0(n3929), .B1(
        image_data[482]), .Y(n3930) );
  AOI22XL U4968 ( .A0(n3896), .A1(image_data[127]), .B0(n3897), .B1(
        image_data[255]), .Y(n4392) );
  AOI22XL U4969 ( .A0(n4763), .A1(image_data[111]), .B0(n3888), .B1(
        image_data[239]), .Y(n4388) );
  AOI22XL U4970 ( .A0(n4721), .A1(image_data[119]), .B0(n3879), .B1(
        image_data[247]), .Y(n4384) );
  AOI22XL U4971 ( .A0(n4714), .A1(image_data[103]), .B0(n3869), .B1(
        image_data[231]), .Y(n4380) );
  AOI22XL U4972 ( .A0(n4702), .A1(image_data[351]), .B0(n3894), .B1(
        image_data[479]), .Y(n4374) );
  AOI22XL U4973 ( .A0(n4763), .A1(image_data[367]), .B0(n3888), .B1(
        image_data[495]), .Y(n4368) );
  AOI22XL U4974 ( .A0(n4721), .A1(image_data[375]), .B0(n3879), .B1(
        image_data[503]), .Y(n4364) );
  AND2XL U4975 ( .A(IROM_A[4]), .B(n4535), .Y(n3404) );
  NAND2XL U4976 ( .A(IROM_A[0]), .B(IROM_A[1]), .Y(n4555) );
  AOI22XL U4977 ( .A0(n3887), .A1(image_data[305]), .B0(n3936), .B1(
        image_data[433]), .Y(n4924) );
  AOI22XL U4978 ( .A0(n3884), .A1(image_data[273]), .B0(n3934), .B1(
        image_data[401]), .Y(n4926) );
  AOI22XL U4979 ( .A0(n3935), .A1(image_data[369]), .B0(n3888), .B1(
        image_data[497]), .Y(n4923) );
  AOI22XL U4980 ( .A0(n3885), .A1(image_data[337]), .B0(n3886), .B1(
        image_data[465]), .Y(n4925) );
  NAND4XL U4981 ( .A(n4942), .B(n4941), .C(n4940), .D(n4939), .Y(n4958) );
  AOI22XL U4982 ( .A0(n3928), .A1(image_data[33]), .B0(n3929), .B1(
        image_data[161]), .Y(n4940) );
  AOI22XL U4983 ( .A0(n3897), .A1(image_data[1]), .B0(n3896), .B1(
        image_data[129]), .Y(n4942) );
  AOI22XL U4984 ( .A0(n3893), .A1(image_data[97]), .B0(n3894), .B1(
        image_data[225]), .Y(n4939) );
  NAND4XL U4985 ( .A(n4954), .B(n4953), .C(n4952), .D(n4951), .Y(n4955) );
  AOI22XL U4986 ( .A0(n3875), .A1(image_data[89]), .B0(n3876), .B1(
        image_data[217]), .Y(n4953) );
  AOI22XL U4987 ( .A0(n3878), .A1(image_data[121]), .B0(n3879), .B1(
        image_data[249]), .Y(n4951) );
  AOI22XL U4988 ( .A0(n3877), .A1(image_data[57]), .B0(n3949), .B1(
        image_data[185]), .Y(n4952) );
  NAND4XL U4989 ( .A(n4946), .B(n4945), .C(n4944), .D(n4943), .Y(n4957) );
  AOI22XL U4990 ( .A0(n3885), .A1(image_data[81]), .B0(n3886), .B1(
        image_data[209]), .Y(n4945) );
  AOI22XL U4991 ( .A0(n3935), .A1(image_data[113]), .B0(n3888), .B1(
        image_data[241]), .Y(n4943) );
  AOI22XL U4992 ( .A0(n3884), .A1(image_data[17]), .B0(n3934), .B1(
        image_data[145]), .Y(n4946) );
  NAND4XL U4993 ( .A(n4950), .B(n4949), .C(n4948), .D(n4947), .Y(n4956) );
  AOI22XL U4994 ( .A0(n3866), .A1(image_data[73]), .B0(n3867), .B1(
        image_data[201]), .Y(n4949) );
  AOI22XL U4995 ( .A0(n3865), .A1(image_data[9]), .B0(n3941), .B1(
        image_data[137]), .Y(n4950) );
  AOI22XL U4996 ( .A0(n3868), .A1(image_data[105]), .B0(n3869), .B1(
        image_data[233]), .Y(n4947) );
  NAND4XL U4997 ( .A(n4922), .B(n4921), .C(n4920), .D(n4919), .Y(n4938) );
  AOI22XL U4998 ( .A0(n4702), .A1(image_data[353]), .B0(n3894), .B1(
        image_data[481]), .Y(n4919) );
  AOI22XL U4999 ( .A0(n3928), .A1(image_data[289]), .B0(n3929), .B1(
        image_data[417]), .Y(n4920) );
  AOI22XL U5000 ( .A0(n3897), .A1(image_data[257]), .B0(n3896), .B1(
        image_data[385]), .Y(n4922) );
  NAND4XL U5001 ( .A(n4934), .B(n4933), .C(n4932), .D(n4931), .Y(n4935) );
  AOI22XL U5002 ( .A0(n3875), .A1(image_data[345]), .B0(n3876), .B1(
        image_data[473]), .Y(n4933) );
  AOI22XL U5003 ( .A0(n3877), .A1(image_data[313]), .B0(n3949), .B1(
        image_data[441]), .Y(n4932) );
  AOI22XL U5004 ( .A0(n3874), .A1(image_data[281]), .B0(n3948), .B1(
        image_data[409]), .Y(n4934) );
  NAND4XL U5005 ( .A(n4930), .B(n4929), .C(n4928), .D(n4927), .Y(n4936) );
  AOI22XL U5006 ( .A0(n3866), .A1(image_data[329]), .B0(n3867), .B1(
        image_data[457]), .Y(n4929) );
  AOI22XL U5007 ( .A0(n3865), .A1(image_data[265]), .B0(n3941), .B1(
        image_data[393]), .Y(n4930) );
  AOI22XL U5008 ( .A0(n3942), .A1(image_data[297]), .B0(n3943), .B1(
        image_data[425]), .Y(n4928) );
  AOI22XL U5009 ( .A0(n3884), .A1(image_data[329]), .B0(n3934), .B1(
        image_data[457]), .Y(n4648) );
  AOI22XL U5010 ( .A0(n3887), .A1(image_data[361]), .B0(n3936), .B1(
        image_data[489]), .Y(n4646) );
  AOI22XL U5011 ( .A0(n3888), .A1(image_data[297]), .B0(n4763), .B1(
        image_data[425]), .Y(n4647) );
  AOI22XL U5012 ( .A0(n3886), .A1(image_data[265]), .B0(n3885), .B1(
        image_data[393]), .Y(n4649) );
  NAND4XL U5013 ( .A(n4674), .B(n4673), .C(n4672), .D(n4671), .Y(n4675) );
  AOI22XL U5014 ( .A0(n4670), .A1(image_data[57]), .B0(n3896), .B1(
        image_data[185]), .Y(n4672) );
  AOI22XL U5015 ( .A0(n3928), .A1(image_data[89]), .B0(n3929), .B1(
        image_data[217]), .Y(n4673) );
  AOI22XL U5016 ( .A0(n3894), .A1(image_data[25]), .B0(n3893), .B1(
        image_data[153]), .Y(n4674) );
  NAND4XL U5017 ( .A(n4665), .B(n4664), .C(n4663), .D(n4662), .Y(n4677) );
  AOI22XL U5018 ( .A0(n3876), .A1(image_data[17]), .B0(n3875), .B1(
        image_data[145]), .Y(n4665) );
  AOI22XL U5019 ( .A0(n3877), .A1(image_data[113]), .B0(n3949), .B1(
        image_data[241]), .Y(n4662) );
  AOI22XL U5020 ( .A0(n3874), .A1(image_data[81]), .B0(n3948), .B1(
        image_data[209]), .Y(n4664) );
  NAND4XL U5021 ( .A(n4661), .B(n4660), .C(n4659), .D(n4658), .Y(n4678) );
  AOI22XL U5022 ( .A0(n3867), .A1(image_data[1]), .B0(n3866), .B1(
        image_data[129]), .Y(n4661) );
  AOI22XL U5023 ( .A0(n3865), .A1(image_data[65]), .B0(n3941), .B1(
        image_data[193]), .Y(n4660) );
  AOI22XL U5024 ( .A0(n3942), .A1(image_data[97]), .B0(n3943), .B1(
        image_data[225]), .Y(n4658) );
  NAND4XL U5025 ( .A(n4669), .B(n4668), .C(n4667), .D(n4666), .Y(n4676) );
  AOI22XL U5026 ( .A0(n3886), .A1(image_data[9]), .B0(n3885), .B1(
        image_data[137]), .Y(n4669) );
  AOI22XL U5027 ( .A0(n3888), .A1(image_data[41]), .B0(n4763), .B1(
        image_data[169]), .Y(n4667) );
  AOI22XL U5028 ( .A0(n3887), .A1(image_data[105]), .B0(n3936), .B1(
        image_data[233]), .Y(n4666) );
  NAND4XL U5029 ( .A(n4653), .B(n4652), .C(n4651), .D(n4650), .Y(n4654) );
  AOI22XL U5030 ( .A0(n3897), .A1(image_data[313]), .B0(n4768), .B1(
        image_data[441]), .Y(n4651) );
  AOI22XL U5031 ( .A0(n3928), .A1(image_data[345]), .B0(n3929), .B1(
        image_data[473]), .Y(n4652) );
  AOI22XL U5032 ( .A0(n3894), .A1(image_data[281]), .B0(n3893), .B1(
        image_data[409]), .Y(n4653) );
  NAND4XL U5033 ( .A(n4645), .B(n4644), .C(n4643), .D(n4642), .Y(n4656) );
  AOI22XL U5034 ( .A0(n3876), .A1(image_data[273]), .B0(n3875), .B1(
        image_data[401]), .Y(n4645) );
  AOI22XL U5035 ( .A0(n3877), .A1(image_data[369]), .B0(n3949), .B1(
        image_data[497]), .Y(n4642) );
  AOI22XL U5036 ( .A0(n3874), .A1(image_data[337]), .B0(n3948), .B1(
        image_data[465]), .Y(n4644) );
  NAND4XL U5037 ( .A(n4641), .B(n4640), .C(n4639), .D(n4638), .Y(n4657) );
  AOI22XL U5038 ( .A0(n3867), .A1(image_data[257]), .B0(n3866), .B1(
        image_data[385]), .Y(n4641) );
  AOI22XL U5039 ( .A0(n4753), .A1(image_data[321]), .B0(n3941), .B1(
        image_data[449]), .Y(n4640) );
  AOI22XL U5040 ( .A0(n4754), .A1(image_data[353]), .B0(n3943), .B1(
        image_data[481]), .Y(n4638) );
  AOI22XL U5041 ( .A0(n4721), .A1(image_data[376]), .B0(n3879), .B1(
        image_data[504]), .Y(n4889) );
  AOI22XL U5042 ( .A0(n3874), .A1(image_data[280]), .B0(n3948), .B1(
        image_data[408]), .Y(n4892) );
  AOI22XL U5043 ( .A0(n3877), .A1(image_data[312]), .B0(n3949), .B1(
        image_data[440]), .Y(n4890) );
  AOI22XL U5044 ( .A0(n3875), .A1(image_data[344]), .B0(n3876), .B1(
        image_data[472]), .Y(n4891) );
  NAND4XL U5045 ( .A(n4904), .B(n4903), .C(n4902), .D(n4901), .Y(n4915) );
  AOI22XL U5046 ( .A0(n3885), .A1(image_data[80]), .B0(n3886), .B1(
        image_data[208]), .Y(n4903) );
  AOI22XL U5047 ( .A0(n3884), .A1(image_data[16]), .B0(n3934), .B1(
        image_data[144]), .Y(n4904) );
  AOI22XL U5048 ( .A0(n3887), .A1(image_data[48]), .B0(n3936), .B1(
        image_data[176]), .Y(n4902) );
  NAND4XL U5049 ( .A(n4900), .B(n4899), .C(n4898), .D(n4897), .Y(n4916) );
  AOI22XL U5050 ( .A0(n3928), .A1(image_data[32]), .B0(n3929), .B1(
        image_data[160]), .Y(n4898) );
  AOI22XL U5051 ( .A0(n3897), .A1(image_data[0]), .B0(n3896), .B1(
        image_data[128]), .Y(n4900) );
  AOI22XL U5052 ( .A0(n4702), .A1(image_data[96]), .B0(n3894), .B1(
        image_data[224]), .Y(n4897) );
  NAND4XL U5053 ( .A(n4908), .B(n4907), .C(n4906), .D(n4905), .Y(n4914) );
  AOI22XL U5054 ( .A0(n3865), .A1(image_data[8]), .B0(n3941), .B1(
        image_data[136]), .Y(n4908) );
  AOI22XL U5055 ( .A0(n3866), .A1(image_data[72]), .B0(n3867), .B1(
        image_data[200]), .Y(n4907) );
  AOI22XL U5056 ( .A0(n3942), .A1(image_data[40]), .B0(n3943), .B1(
        image_data[168]), .Y(n4906) );
  NAND4XL U5057 ( .A(n4912), .B(n4911), .C(n4910), .D(n4909), .Y(n4913) );
  AOI22XL U5058 ( .A0(n3875), .A1(image_data[88]), .B0(n3876), .B1(
        image_data[216]), .Y(n4911) );
  AOI22XL U5059 ( .A0(n3877), .A1(image_data[56]), .B0(n3949), .B1(
        image_data[184]), .Y(n4910) );
  AOI22XL U5060 ( .A0(n3874), .A1(image_data[24]), .B0(n3948), .B1(
        image_data[152]), .Y(n4912) );
  NAND4XL U5061 ( .A(n4884), .B(n4883), .C(n4882), .D(n4881), .Y(n4895) );
  AOI22XL U5062 ( .A0(n3885), .A1(image_data[336]), .B0(n3886), .B1(
        image_data[464]), .Y(n4883) );
  AOI22XL U5063 ( .A0(n3884), .A1(image_data[272]), .B0(n3934), .B1(
        image_data[400]), .Y(n4884) );
  AOI22XL U5064 ( .A0(n3887), .A1(image_data[304]), .B0(n3936), .B1(
        image_data[432]), .Y(n4882) );
  NAND4XL U5065 ( .A(n4880), .B(n4879), .C(n4878), .D(n4877), .Y(n4896) );
  AOI22XL U5066 ( .A0(n3928), .A1(image_data[288]), .B0(n3929), .B1(
        image_data[416]), .Y(n4878) );
  AOI22XL U5067 ( .A0(n3897), .A1(image_data[256]), .B0(n3896), .B1(
        image_data[384]), .Y(n4880) );
  AOI22XL U5068 ( .A0(n4702), .A1(image_data[352]), .B0(n3894), .B1(
        image_data[480]), .Y(n4877) );
  NAND4XL U5069 ( .A(n4888), .B(n4887), .C(n4886), .D(n4885), .Y(n4894) );
  AOI22XL U5070 ( .A0(n3865), .A1(image_data[264]), .B0(n3941), .B1(
        image_data[392]), .Y(n4888) );
  AOI22XL U5071 ( .A0(n3866), .A1(image_data[328]), .B0(n3867), .B1(
        image_data[456]), .Y(n4887) );
  AOI22XL U5072 ( .A0(n3942), .A1(image_data[296]), .B0(n3943), .B1(
        image_data[424]), .Y(n4886) );
  AOI22XL U5073 ( .A0(n3884), .A1(image_data[328]), .B0(n3934), .B1(
        image_data[456]), .Y(n4743) );
  AOI22XL U5074 ( .A0(n3887), .A1(image_data[360]), .B0(n3936), .B1(
        image_data[488]), .Y(n4741) );
  AOI22XL U5075 ( .A0(n3888), .A1(image_data[296]), .B0(n4763), .B1(
        image_data[424]), .Y(n4742) );
  AOI22XL U5076 ( .A0(n3886), .A1(image_data[264]), .B0(n3885), .B1(
        image_data[392]), .Y(n4744) );
  NAND4XL U5077 ( .A(n4772), .B(n4771), .C(n4770), .D(n4769), .Y(n4773) );
  AOI22XL U5078 ( .A0(n3897), .A1(image_data[56]), .B0(n4768), .B1(
        image_data[184]), .Y(n4770) );
  AOI22XL U5079 ( .A0(n3928), .A1(image_data[88]), .B0(n3929), .B1(
        image_data[216]), .Y(n4771) );
  AOI22XL U5080 ( .A0(n3894), .A1(image_data[24]), .B0(n3893), .B1(
        image_data[152]), .Y(n4772) );
  NAND4XL U5081 ( .A(n4762), .B(n4761), .C(n4760), .D(n4759), .Y(n4775) );
  AOI22XL U5082 ( .A0(n3876), .A1(image_data[16]), .B0(n3875), .B1(
        image_data[144]), .Y(n4762) );
  AOI22XL U5083 ( .A0(n3877), .A1(image_data[112]), .B0(n3949), .B1(
        image_data[240]), .Y(n4759) );
  AOI22XL U5084 ( .A0(n3874), .A1(image_data[80]), .B0(n3948), .B1(
        image_data[208]), .Y(n4761) );
  NAND4XL U5085 ( .A(n4758), .B(n4757), .C(n4756), .D(n4755), .Y(n4776) );
  AOI22XL U5086 ( .A0(n4753), .A1(image_data[64]), .B0(n3941), .B1(
        image_data[192]), .Y(n4757) );
  AOI22XL U5087 ( .A0(n3867), .A1(image_data[0]), .B0(n3866), .B1(
        image_data[128]), .Y(n4758) );
  AOI22XL U5088 ( .A0(n4754), .A1(image_data[96]), .B0(n3943), .B1(
        image_data[224]), .Y(n4755) );
  NAND4XL U5089 ( .A(n4767), .B(n4766), .C(n4765), .D(n4764), .Y(n4774) );
  AOI22XL U5090 ( .A0(n3886), .A1(image_data[8]), .B0(n3885), .B1(
        image_data[136]), .Y(n4767) );
  AOI22XL U5091 ( .A0(n3888), .A1(image_data[40]), .B0(n4763), .B1(
        image_data[168]), .Y(n4765) );
  AOI22XL U5092 ( .A0(n3887), .A1(image_data[104]), .B0(n3936), .B1(
        image_data[232]), .Y(n4764) );
  NAND4XL U5093 ( .A(n4740), .B(n4739), .C(n4738), .D(n4737), .Y(n4751) );
  AOI22XL U5094 ( .A0(n3876), .A1(image_data[272]), .B0(n3875), .B1(
        image_data[400]), .Y(n4740) );
  AOI22XL U5095 ( .A0(n3877), .A1(image_data[368]), .B0(n3949), .B1(
        image_data[496]), .Y(n4737) );
  AOI22XL U5096 ( .A0(n3874), .A1(image_data[336]), .B0(n3948), .B1(
        image_data[464]), .Y(n4739) );
  NAND4XL U5097 ( .A(n4748), .B(n4747), .C(n4746), .D(n4745), .Y(n4749) );
  AOI22XL U5098 ( .A0(n4681), .A1(image_data[376]), .B0(n3364), .B1(
        image_data[504]), .Y(n4745) );
  AOI22XL U5099 ( .A0(n3897), .A1(image_data[312]), .B0(n4768), .B1(
        image_data[440]), .Y(n4746) );
  AOI22XL U5100 ( .A0(n3928), .A1(image_data[344]), .B0(n3929), .B1(
        image_data[472]), .Y(n4747) );
  NAND4XL U5101 ( .A(n4736), .B(n4735), .C(n4734), .D(n4733), .Y(n4752) );
  AOI22XL U5102 ( .A0(n3865), .A1(image_data[320]), .B0(n3941), .B1(
        image_data[448]), .Y(n4735) );
  AOI22XL U5103 ( .A0(n3867), .A1(image_data[256]), .B0(n3866), .B1(
        image_data[384]), .Y(n4736) );
  AOI22XL U5104 ( .A0(n4754), .A1(image_data[352]), .B0(n3943), .B1(
        image_data[480]), .Y(n4733) );
  OAI2BB1XL U5105 ( .A0N(n5262), .A1N(n5261), .B0(n5260), .Y(n6116) );
  NAND4XL U5106 ( .A(n6043), .B(n6042), .C(n6041), .D(n6040), .Y(n6049) );
  AOI22XL U5107 ( .A0(n6468), .A1(image_data[264]), .B0(n6467), .B1(
        image_data[392]), .Y(n6043) );
  AOI22XL U5108 ( .A0(n6470), .A1(image_data[328]), .B0(n6469), .B1(
        image_data[456]), .Y(n6042) );
  AOI22XL U5109 ( .A0(n6472), .A1(image_data[296]), .B0(n6471), .B1(
        image_data[424]), .Y(n6041) );
  NAND4XL U5110 ( .A(n6047), .B(n6046), .C(n6045), .D(n6044), .Y(n6048) );
  AOI22XL U5111 ( .A0(n6480), .A1(image_data[280]), .B0(n6479), .B1(
        image_data[408]), .Y(n6047) );
  AOI22XL U5112 ( .A0(n6482), .A1(image_data[344]), .B0(n6481), .B1(
        image_data[472]), .Y(n6046) );
  AOI22XL U5113 ( .A0(n6484), .A1(image_data[312]), .B0(n6483), .B1(
        image_data[440]), .Y(n6045) );
  NAND4XL U5114 ( .A(n6035), .B(n6034), .C(n6033), .D(n6032), .Y(n6051) );
  AOI22XL U5115 ( .A0(n6444), .A1(image_data[256]), .B0(n6443), .B1(
        image_data[384]), .Y(n6035) );
  AOI22XL U5116 ( .A0(n6446), .A1(image_data[320]), .B0(n6445), .B1(
        image_data[448]), .Y(n6034) );
  AOI22XL U5117 ( .A0(n6448), .A1(image_data[288]), .B0(n6447), .B1(
        image_data[416]), .Y(n6033) );
  NAND4XL U5118 ( .A(n6039), .B(n6038), .C(n6037), .D(n6036), .Y(n6050) );
  AOI22XL U5119 ( .A0(n6456), .A1(image_data[272]), .B0(n6455), .B1(
        image_data[400]), .Y(n6039) );
  AOI22XL U5120 ( .A0(n6460), .A1(image_data[304]), .B0(n6459), .B1(
        image_data[432]), .Y(n6037) );
  AOI22XL U5121 ( .A0(n6462), .A1(image_data[368]), .B0(n6461), .B1(
        image_data[496]), .Y(n6036) );
  NOR4XL U5122 ( .A(n6113), .B(n6112), .C(n6111), .D(n6110), .Y(n6114) );
  NAND4XL U5123 ( .A(n6101), .B(n6100), .C(n6099), .D(n6098), .Y(n6112) );
  NAND4XL U5124 ( .A(n6097), .B(n6096), .C(n6095), .D(n6094), .Y(n6113) );
  NAND4XL U5125 ( .A(n6109), .B(n6108), .C(n6107), .D(n6106), .Y(n6110) );
  NOR4XL U5126 ( .A(n6093), .B(n6092), .C(n6091), .D(n6090), .Y(n6115) );
  NAND4XL U5127 ( .A(n6081), .B(n6080), .C(n6079), .D(n6078), .Y(n6092) );
  NAND4XL U5128 ( .A(n6077), .B(n6076), .C(n6075), .D(n6074), .Y(n6093) );
  NAND4XL U5129 ( .A(n6089), .B(n6088), .C(n6087), .D(n6086), .Y(n6090) );
  NOR4XL U5130 ( .A(n6071), .B(n6070), .C(n6069), .D(n6068), .Y(n6072) );
  NAND4XL U5131 ( .A(n6059), .B(n6058), .C(n6057), .D(n6056), .Y(n6070) );
  NAND4XL U5132 ( .A(n6055), .B(n6054), .C(n6053), .D(n6052), .Y(n6071) );
  NAND4XL U5133 ( .A(n6067), .B(n6066), .C(n6065), .D(n6064), .Y(n6068) );
  NAND4XL U5134 ( .A(n4863), .B(n4862), .C(n4861), .D(n4860), .Y(n4864) );
  AOI22XL U5135 ( .A0(n4702), .A1(image_data[89]), .B0(n3894), .B1(
        image_data[217]), .Y(n4862) );
  AOI22XL U5136 ( .A0(n3896), .A1(image_data[121]), .B0(n3897), .B1(
        image_data[249]), .Y(n4860) );
  AOI22XL U5137 ( .A0(n3928), .A1(image_data[25]), .B0(n3929), .B1(
        image_data[153]), .Y(n4863) );
  NAND4XL U5138 ( .A(n4859), .B(n4858), .C(n4857), .D(n4856), .Y(n4865) );
  AOI22XL U5139 ( .A0(n4707), .A1(image_data[73]), .B0(n3886), .B1(
        image_data[201]), .Y(n4858) );
  AOI22XL U5140 ( .A0(n3935), .A1(image_data[105]), .B0(n3888), .B1(
        image_data[233]), .Y(n4856) );
  AOI22XL U5141 ( .A0(n3884), .A1(image_data[9]), .B0(n3934), .B1(
        image_data[137]), .Y(n4859) );
  NAND4XL U5142 ( .A(n4855), .B(n4854), .C(n4853), .D(n4852), .Y(n4866) );
  AOI22XL U5143 ( .A0(n4719), .A1(image_data[81]), .B0(n3876), .B1(
        image_data[209]), .Y(n4854) );
  AOI22XL U5144 ( .A0(n3877), .A1(image_data[49]), .B0(n3949), .B1(
        image_data[177]), .Y(n4853) );
  AOI22XL U5145 ( .A0(n3874), .A1(image_data[17]), .B0(n3948), .B1(
        image_data[145]), .Y(n4855) );
  NAND4XL U5146 ( .A(n4851), .B(n4850), .C(n4849), .D(n4848), .Y(n4867) );
  AOI22XL U5147 ( .A0(n3866), .A1(image_data[65]), .B0(n3867), .B1(
        image_data[193]), .Y(n4850) );
  AOI22XL U5148 ( .A0(n3865), .A1(image_data[1]), .B0(n3941), .B1(
        image_data[129]), .Y(n4851) );
  AOI22XL U5149 ( .A0(n3942), .A1(image_data[33]), .B0(n3943), .B1(
        image_data[161]), .Y(n4849) );
  NAND4XL U5150 ( .A(n4843), .B(n4842), .C(n4841), .D(n4840), .Y(n4844) );
  AOI22XL U5151 ( .A0(n3896), .A1(image_data[377]), .B0(n3897), .B1(
        image_data[505]), .Y(n4840) );
  AOI22XL U5152 ( .A0(n3928), .A1(image_data[281]), .B0(n3929), .B1(
        image_data[409]), .Y(n4843) );
  AOI22XL U5153 ( .A0(n3893), .A1(image_data[345]), .B0(n3894), .B1(
        image_data[473]), .Y(n4842) );
  NAND4XL U5154 ( .A(n4839), .B(n4838), .C(n4837), .D(n4836), .Y(n4845) );
  AOI22XL U5155 ( .A0(n4707), .A1(image_data[329]), .B0(n3886), .B1(
        image_data[457]), .Y(n4838) );
  AOI22XL U5156 ( .A0(n3935), .A1(image_data[361]), .B0(n3888), .B1(
        image_data[489]), .Y(n4836) );
  AOI22XL U5157 ( .A0(n3884), .A1(image_data[265]), .B0(n3934), .B1(
        image_data[393]), .Y(n4839) );
  NAND4XL U5158 ( .A(n4835), .B(n4834), .C(n4833), .D(n4832), .Y(n4846) );
  AOI22XL U5159 ( .A0(n3875), .A1(image_data[337]), .B0(n3876), .B1(
        image_data[465]), .Y(n4834) );
  AOI22XL U5160 ( .A0(n3877), .A1(image_data[305]), .B0(n3949), .B1(
        image_data[433]), .Y(n4833) );
  AOI22XL U5161 ( .A0(n3874), .A1(image_data[273]), .B0(n3948), .B1(
        image_data[401]), .Y(n4835) );
  NAND4XL U5162 ( .A(n4831), .B(n4830), .C(n4829), .D(n4828), .Y(n4847) );
  AOI22XL U5163 ( .A0(n3866), .A1(image_data[321]), .B0(n3867), .B1(
        image_data[449]), .Y(n4830) );
  AOI22XL U5164 ( .A0(n3865), .A1(image_data[257]), .B0(n3941), .B1(
        image_data[385]), .Y(n4831) );
  AOI22XL U5165 ( .A0(n3942), .A1(image_data[289]), .B0(n3943), .B1(
        image_data[417]), .Y(n4829) );
  AOI22XL U5166 ( .A0(n3884), .A1(image_data[337]), .B0(n3934), .B1(
        image_data[465]), .Y(n4688) );
  AOI22XL U5167 ( .A0(n3888), .A1(image_data[305]), .B0(n3935), .B1(
        image_data[433]), .Y(n4687) );
  AOI22XL U5168 ( .A0(n3887), .A1(image_data[369]), .B0(n3936), .B1(
        image_data[497]), .Y(n4686) );
  AOI22XL U5169 ( .A0(n3886), .A1(image_data[273]), .B0(n3885), .B1(
        image_data[401]), .Y(n4689) );
  NAND4XL U5170 ( .A(n4706), .B(n4705), .C(n4704), .D(n4703), .Y(n4730) );
  AOI22XL U5171 ( .A0(n3894), .A1(image_data[33]), .B0(n4702), .B1(
        image_data[161]), .Y(n4704) );
  AOI22XL U5172 ( .A0(n3897), .A1(image_data[65]), .B0(n3896), .B1(
        image_data[193]), .Y(n4705) );
  AOI22XL U5173 ( .A0(n3928), .A1(image_data[97]), .B0(n3929), .B1(
        image_data[225]), .Y(n4703) );
  NAND4XL U5174 ( .A(n4726), .B(n4725), .C(n4724), .D(n4723), .Y(n4727) );
  AOI22XL U5175 ( .A0(n3876), .A1(image_data[25]), .B0(n4719), .B1(
        image_data[153]), .Y(n4726) );
  AOI22XL U5176 ( .A0(n3879), .A1(image_data[57]), .B0(n4721), .B1(
        image_data[185]), .Y(n4724) );
  AOI22XL U5177 ( .A0(n4722), .A1(image_data[121]), .B0(n3949), .B1(
        image_data[249]), .Y(n4723) );
  NAND4XL U5178 ( .A(n4718), .B(n4717), .C(n4716), .D(n4715), .Y(n4728) );
  AOI22XL U5179 ( .A0(n3867), .A1(image_data[9]), .B0(n4713), .B1(
        image_data[137]), .Y(n4718) );
  AOI22XL U5180 ( .A0(n3869), .A1(image_data[41]), .B0(n4714), .B1(
        image_data[169]), .Y(n4716) );
  AOI22XL U5181 ( .A0(n3865), .A1(image_data[73]), .B0(n3941), .B1(
        image_data[201]), .Y(n4717) );
  NAND4XL U5182 ( .A(n4712), .B(n4711), .C(n4710), .D(n4709), .Y(n4729) );
  AOI22XL U5183 ( .A0(n3886), .A1(image_data[17]), .B0(n4707), .B1(
        image_data[145]), .Y(n4712) );
  AOI22XL U5184 ( .A0(n3887), .A1(image_data[113]), .B0(n3936), .B1(
        image_data[241]), .Y(n4709) );
  AOI22XL U5185 ( .A0(n3888), .A1(image_data[49]), .B0(n3935), .B1(
        image_data[177]), .Y(n4710) );
  NAND4XL U5186 ( .A(n4697), .B(n4696), .C(n4695), .D(n4694), .Y(n4698) );
  AOI22XL U5187 ( .A0(n3876), .A1(image_data[281]), .B0(n4719), .B1(
        image_data[409]), .Y(n4697) );
  AOI22XL U5188 ( .A0(n3879), .A1(image_data[313]), .B0(n4721), .B1(
        image_data[441]), .Y(n4695) );
  AOI22XL U5189 ( .A0(n4722), .A1(image_data[377]), .B0(n3949), .B1(
        image_data[505]), .Y(n4694) );
  NAND4XL U5190 ( .A(n4693), .B(n4692), .C(n4691), .D(n4690), .Y(n4699) );
  AOI22XL U5191 ( .A0(n3867), .A1(image_data[265]), .B0(n4713), .B1(
        image_data[393]), .Y(n4693) );
  AOI22XL U5192 ( .A0(n3869), .A1(image_data[297]), .B0(n4714), .B1(
        image_data[425]), .Y(n4691) );
  AOI22XL U5193 ( .A0(n3865), .A1(image_data[329]), .B0(n3941), .B1(
        image_data[457]), .Y(n4692) );
  NAND4XL U5194 ( .A(n4685), .B(n4684), .C(n4683), .D(n4682), .Y(n4701) );
  AOI22XL U5195 ( .A0(n3364), .A1(image_data[257]), .B0(n4681), .B1(
        image_data[385]), .Y(n4685) );
  AOI22XL U5196 ( .A0(n3897), .A1(image_data[321]), .B0(n3896), .B1(
        image_data[449]), .Y(n4684) );
  AOI22XL U5197 ( .A0(n3928), .A1(image_data[353]), .B0(n3929), .B1(
        image_data[481]), .Y(n4682) );
  AOI22XL U5198 ( .A0(n6486), .A1(image_data[123]), .B0(n6485), .B1(
        image_data[251]), .Y(n6209) );
  AOI22XL U5199 ( .A0(n6484), .A1(image_data[59]), .B0(n6483), .B1(
        image_data[187]), .Y(n6210) );
  AOI22XL U5200 ( .A0(n6482), .A1(image_data[91]), .B0(n6481), .B1(
        image_data[219]), .Y(n6211) );
  AOI22XL U5201 ( .A0(n6480), .A1(image_data[27]), .B0(n6479), .B1(
        image_data[155]), .Y(n6212) );
  AOI22XL U5202 ( .A0(n6450), .A1(image_data[99]), .B0(n6449), .B1(
        image_data[227]), .Y(n6197) );
  AOI22XL U5203 ( .A0(n6448), .A1(image_data[35]), .B0(n6447), .B1(
        image_data[163]), .Y(n6198) );
  AOI22XL U5204 ( .A0(n6446), .A1(image_data[67]), .B0(n6445), .B1(
        image_data[195]), .Y(n6199) );
  AOI22XL U5205 ( .A0(n6444), .A1(image_data[3]), .B0(n6443), .B1(
        image_data[131]), .Y(n6200) );
  AOI22XL U5206 ( .A0(n6462), .A1(image_data[115]), .B0(n6461), .B1(
        image_data[243]), .Y(n6201) );
  AOI22XL U5207 ( .A0(n6460), .A1(image_data[51]), .B0(n6459), .B1(
        image_data[179]), .Y(n6202) );
  AOI22XL U5208 ( .A0(n6458), .A1(image_data[83]), .B0(n6457), .B1(
        image_data[211]), .Y(n6203) );
  AOI22XL U5209 ( .A0(n6456), .A1(image_data[19]), .B0(n6455), .B1(
        image_data[147]), .Y(n6204) );
  NAND4XL U5210 ( .A(n6208), .B(n6207), .C(n6206), .D(n6205), .Y(n6214) );
  AOI22XL U5211 ( .A0(n6468), .A1(image_data[11]), .B0(n6467), .B1(
        image_data[139]), .Y(n6208) );
  AOI22XL U5212 ( .A0(n6470), .A1(image_data[75]), .B0(n6469), .B1(
        image_data[203]), .Y(n6207) );
  AOI22XL U5213 ( .A0(n6472), .A1(image_data[43]), .B0(n6471), .B1(
        image_data[171]), .Y(n6206) );
  AOI22XL U5214 ( .A0(n6486), .A1(image_data[379]), .B0(n6485), .B1(
        image_data[507]), .Y(n6189) );
  AOI22XL U5215 ( .A0(n6484), .A1(image_data[315]), .B0(n6483), .B1(
        image_data[443]), .Y(n6190) );
  AOI22XL U5216 ( .A0(n6482), .A1(image_data[347]), .B0(n6481), .B1(
        image_data[475]), .Y(n6191) );
  AOI22XL U5217 ( .A0(n6480), .A1(image_data[283]), .B0(n6479), .B1(
        image_data[411]), .Y(n6192) );
  AOI22XL U5218 ( .A0(n6462), .A1(image_data[371]), .B0(n6461), .B1(
        image_data[499]), .Y(n6181) );
  AOI22XL U5219 ( .A0(n6460), .A1(image_data[307]), .B0(n6459), .B1(
        image_data[435]), .Y(n6182) );
  AOI22XL U5220 ( .A0(n6458), .A1(image_data[339]), .B0(n6457), .B1(
        image_data[467]), .Y(n6183) );
  AOI22XL U5221 ( .A0(n6456), .A1(image_data[275]), .B0(n6455), .B1(
        image_data[403]), .Y(n6184) );
  AOI22XL U5222 ( .A0(n6450), .A1(image_data[355]), .B0(n6449), .B1(
        image_data[483]), .Y(n6177) );
  AOI22XL U5223 ( .A0(n6448), .A1(image_data[291]), .B0(n6447), .B1(
        image_data[419]), .Y(n6178) );
  AOI22XL U5224 ( .A0(n6446), .A1(image_data[323]), .B0(n6445), .B1(
        image_data[451]), .Y(n6179) );
  AOI22XL U5225 ( .A0(n6444), .A1(image_data[259]), .B0(n6443), .B1(
        image_data[387]), .Y(n6180) );
  NAND4XL U5226 ( .A(n6188), .B(n6187), .C(n6186), .D(n6185), .Y(n6194) );
  AOI22XL U5227 ( .A0(n6468), .A1(image_data[267]), .B0(n6467), .B1(
        image_data[395]), .Y(n6188) );
  AOI22XL U5228 ( .A0(n6470), .A1(image_data[331]), .B0(n6469), .B1(
        image_data[459]), .Y(n6187) );
  AOI22XL U5229 ( .A0(n6472), .A1(image_data[299]), .B0(n6471), .B1(
        image_data[427]), .Y(n6186) );
  AOI22XL U5230 ( .A0(n6534), .A1(image_data[339]), .B0(n6533), .B1(
        image_data[467]), .Y(n6225) );
  AOI22XL U5231 ( .A0(n6538), .A1(image_data[371]), .B0(n6537), .B1(
        image_data[499]), .Y(n6223) );
  AOI22XL U5232 ( .A0(n6536), .A1(image_data[307]), .B0(n6535), .B1(
        image_data[435]), .Y(n6224) );
  AOI22XL U5233 ( .A0(n6532), .A1(image_data[275]), .B0(n6531), .B1(
        image_data[403]), .Y(n6226) );
  NAND4XL U5234 ( .A(n6250), .B(n6249), .C(n6248), .D(n6247), .Y(n6256) );
  AOI22XL U5235 ( .A0(n6544), .A1(image_data[11]), .B0(n6543), .B1(
        image_data[139]), .Y(n6250) );
  AOI22XL U5236 ( .A0(n6546), .A1(image_data[75]), .B0(n6545), .B1(
        image_data[203]), .Y(n6249) );
  AOI22XL U5237 ( .A0(n6548), .A1(image_data[43]), .B0(n6547), .B1(
        image_data[171]), .Y(n6248) );
  NAND4XL U5238 ( .A(n6254), .B(n6253), .C(n6252), .D(n6251), .Y(n6255) );
  AOI22XL U5239 ( .A0(n6556), .A1(image_data[27]), .B0(n6555), .B1(
        image_data[155]), .Y(n6254) );
  AOI22XL U5240 ( .A0(n6558), .A1(image_data[91]), .B0(n6557), .B1(
        image_data[219]), .Y(n6253) );
  AOI22XL U5241 ( .A0(n6560), .A1(image_data[59]), .B0(n6559), .B1(
        image_data[187]), .Y(n6252) );
  NAND4XL U5242 ( .A(n6242), .B(n6241), .C(n6240), .D(n6239), .Y(n6258) );
  AOI22XL U5243 ( .A0(n6520), .A1(image_data[3]), .B0(n6519), .B1(
        image_data[131]), .Y(n6242) );
  AOI22XL U5244 ( .A0(n6522), .A1(image_data[67]), .B0(n6521), .B1(
        image_data[195]), .Y(n6241) );
  AOI22XL U5245 ( .A0(n6524), .A1(image_data[35]), .B0(n6523), .B1(
        image_data[163]), .Y(n6240) );
  NAND4XL U5246 ( .A(n6246), .B(n6245), .C(n6244), .D(n6243), .Y(n6257) );
  AOI22XL U5247 ( .A0(n6532), .A1(image_data[19]), .B0(n6531), .B1(
        image_data[147]), .Y(n6246) );
  AOI22XL U5248 ( .A0(n6536), .A1(image_data[51]), .B0(n6535), .B1(
        image_data[179]), .Y(n6244) );
  AOI22XL U5249 ( .A0(n6538), .A1(image_data[115]), .B0(n6537), .B1(
        image_data[243]), .Y(n6243) );
  NAND4XL U5250 ( .A(n6230), .B(n6229), .C(n6228), .D(n6227), .Y(n6236) );
  AOI22XL U5251 ( .A0(n6544), .A1(image_data[267]), .B0(n6543), .B1(
        image_data[395]), .Y(n6230) );
  AOI22XL U5252 ( .A0(n6546), .A1(image_data[331]), .B0(n6545), .B1(
        image_data[459]), .Y(n6229) );
  AOI22XL U5253 ( .A0(n6548), .A1(image_data[299]), .B0(n6547), .B1(
        image_data[427]), .Y(n6228) );
  NAND4XL U5254 ( .A(n6234), .B(n6233), .C(n6232), .D(n6231), .Y(n6235) );
  AOI22XL U5255 ( .A0(n6556), .A1(image_data[283]), .B0(n6555), .B1(
        image_data[411]), .Y(n6234) );
  AOI22XL U5256 ( .A0(n6558), .A1(image_data[347]), .B0(n6557), .B1(
        image_data[475]), .Y(n6233) );
  AOI22XL U5257 ( .A0(n6560), .A1(image_data[315]), .B0(n6559), .B1(
        image_data[443]), .Y(n6232) );
  NAND4XL U5258 ( .A(n6222), .B(n6221), .C(n6220), .D(n6219), .Y(n6238) );
  AOI22XL U5259 ( .A0(n6520), .A1(image_data[259]), .B0(n6519), .B1(
        image_data[387]), .Y(n6222) );
  AOI22XL U5260 ( .A0(n6522), .A1(image_data[323]), .B0(n6521), .B1(
        image_data[451]), .Y(n6221) );
  AOI22XL U5261 ( .A0(n6524), .A1(image_data[291]), .B0(n6523), .B1(
        image_data[419]), .Y(n6220) );
  NAND4XL U5262 ( .A(n5824), .B(n5823), .C(n5822), .D(n5821), .Y(n5830) );
  AOI22XL U5263 ( .A0(n6468), .A1(image_data[270]), .B0(n6467), .B1(
        image_data[398]), .Y(n5824) );
  AOI22XL U5264 ( .A0(n6470), .A1(image_data[334]), .B0(n6469), .B1(
        image_data[462]), .Y(n5823) );
  AOI22XL U5265 ( .A0(n6472), .A1(image_data[302]), .B0(n6471), .B1(
        image_data[430]), .Y(n5822) );
  NAND4XL U5266 ( .A(n5828), .B(n5827), .C(n5826), .D(n5825), .Y(n5829) );
  AOI22XL U5267 ( .A0(n6480), .A1(image_data[286]), .B0(n6479), .B1(
        image_data[414]), .Y(n5828) );
  AOI22XL U5268 ( .A0(n6482), .A1(image_data[350]), .B0(n6481), .B1(
        image_data[478]), .Y(n5827) );
  AOI22XL U5269 ( .A0(n6484), .A1(image_data[318]), .B0(n6483), .B1(
        image_data[446]), .Y(n5826) );
  NAND4XL U5270 ( .A(n5816), .B(n5815), .C(n5814), .D(n5813), .Y(n5832) );
  AOI22XL U5271 ( .A0(n6444), .A1(image_data[262]), .B0(n6443), .B1(
        image_data[390]), .Y(n5816) );
  AOI22XL U5272 ( .A0(n6446), .A1(image_data[326]), .B0(n6445), .B1(
        image_data[454]), .Y(n5815) );
  AOI22XL U5273 ( .A0(n6448), .A1(image_data[294]), .B0(n6447), .B1(
        image_data[422]), .Y(n5814) );
  NAND4XL U5274 ( .A(n5820), .B(n5819), .C(n5818), .D(n5817), .Y(n5831) );
  AOI22XL U5275 ( .A0(n6456), .A1(image_data[278]), .B0(n6455), .B1(
        image_data[406]), .Y(n5820) );
  AOI22XL U5276 ( .A0(n6460), .A1(image_data[310]), .B0(n6459), .B1(
        image_data[438]), .Y(n5818) );
  AOI22XL U5277 ( .A0(n6462), .A1(image_data[374]), .B0(n6461), .B1(
        image_data[502]), .Y(n5817) );
  NOR4XL U5278 ( .A(n5894), .B(n5893), .C(n5892), .D(n5891), .Y(n5895) );
  NAND4XL U5279 ( .A(n5882), .B(n5881), .C(n5880), .D(n5879), .Y(n5893) );
  NAND4XL U5280 ( .A(n5878), .B(n5877), .C(n5876), .D(n5875), .Y(n5894) );
  NAND4XL U5281 ( .A(n5890), .B(n5889), .C(n5888), .D(n5887), .Y(n5891) );
  NOR4XL U5282 ( .A(n5874), .B(n5873), .C(n5872), .D(n5871), .Y(n5896) );
  NAND4XL U5283 ( .A(n5862), .B(n5861), .C(n5860), .D(n5859), .Y(n5873) );
  NAND4XL U5284 ( .A(n5858), .B(n5857), .C(n5856), .D(n5855), .Y(n5874) );
  NAND4XL U5285 ( .A(n5870), .B(n5869), .C(n5868), .D(n5867), .Y(n5871) );
  NOR4XL U5286 ( .A(n5852), .B(n5851), .C(n5850), .D(n5849), .Y(n5853) );
  NAND4XL U5287 ( .A(n5840), .B(n5839), .C(n5838), .D(n5837), .Y(n5851) );
  NAND4XL U5288 ( .A(n5836), .B(n5835), .C(n5834), .D(n5833), .Y(n5852) );
  NAND4XL U5289 ( .A(n5848), .B(n5847), .C(n5846), .D(n5845), .Y(n5849) );
  NAND4XL U5290 ( .A(n5619), .B(n5618), .C(n5617), .D(n5616), .Y(n5625) );
  AOI22XL U5291 ( .A0(n6468), .A1(image_data[265]), .B0(n6467), .B1(
        image_data[393]), .Y(n5619) );
  AOI22XL U5292 ( .A0(n6470), .A1(image_data[329]), .B0(n6469), .B1(
        image_data[457]), .Y(n5618) );
  AOI22XL U5293 ( .A0(n6472), .A1(image_data[297]), .B0(n6471), .B1(
        image_data[425]), .Y(n5617) );
  NAND4XL U5294 ( .A(n5623), .B(n5622), .C(n5621), .D(n5620), .Y(n5624) );
  AOI22XL U5295 ( .A0(n6480), .A1(image_data[281]), .B0(n6479), .B1(
        image_data[409]), .Y(n5623) );
  AOI22XL U5296 ( .A0(n6482), .A1(image_data[345]), .B0(n6481), .B1(
        image_data[473]), .Y(n5622) );
  AOI22XL U5297 ( .A0(n6484), .A1(image_data[313]), .B0(n6483), .B1(
        image_data[441]), .Y(n5621) );
  NAND4XL U5298 ( .A(n5611), .B(n5610), .C(n5609), .D(n5608), .Y(n5627) );
  AOI22XL U5299 ( .A0(n6444), .A1(image_data[257]), .B0(n6443), .B1(
        image_data[385]), .Y(n5611) );
  AOI22XL U5300 ( .A0(n6446), .A1(image_data[321]), .B0(n6445), .B1(
        image_data[449]), .Y(n5610) );
  AOI22XL U5301 ( .A0(n6448), .A1(image_data[289]), .B0(n6447), .B1(
        image_data[417]), .Y(n5609) );
  NAND4XL U5302 ( .A(n5615), .B(n5614), .C(n5613), .D(n5612), .Y(n5626) );
  AOI22XL U5303 ( .A0(n6456), .A1(image_data[273]), .B0(n6455), .B1(
        image_data[401]), .Y(n5615) );
  AOI22XL U5304 ( .A0(n6460), .A1(image_data[305]), .B0(n6459), .B1(
        image_data[433]), .Y(n5613) );
  AOI22XL U5305 ( .A0(n6462), .A1(image_data[369]), .B0(n6461), .B1(
        image_data[497]), .Y(n5612) );
  NOR4XL U5306 ( .A(n5689), .B(n5688), .C(n5687), .D(n5686), .Y(n5690) );
  NAND4XL U5307 ( .A(n5677), .B(n5676), .C(n5675), .D(n5674), .Y(n5688) );
  NAND4XL U5308 ( .A(n5673), .B(n5672), .C(n5671), .D(n5670), .Y(n5689) );
  NAND4XL U5309 ( .A(n5685), .B(n5684), .C(n5683), .D(n5682), .Y(n5686) );
  NOR4XL U5310 ( .A(n5669), .B(n5668), .C(n5667), .D(n5666), .Y(n5691) );
  NAND4XL U5311 ( .A(n5657), .B(n5656), .C(n5655), .D(n5654), .Y(n5668) );
  NAND4XL U5312 ( .A(n5653), .B(n5652), .C(n5651), .D(n5650), .Y(n5669) );
  NAND4XL U5313 ( .A(n5665), .B(n5664), .C(n5663), .D(n5662), .Y(n5666) );
  NOR4XL U5314 ( .A(n5647), .B(n5646), .C(n5645), .D(n5644), .Y(n5648) );
  NAND4XL U5315 ( .A(n5635), .B(n5634), .C(n5633), .D(n5632), .Y(n5646) );
  NAND4XL U5316 ( .A(n5631), .B(n5630), .C(n5629), .D(n5628), .Y(n5647) );
  NAND4XL U5317 ( .A(n5643), .B(n5642), .C(n5641), .D(n5640), .Y(n5644) );
  AOI22XL U5318 ( .A0(n6526), .A1(image_data[359]), .B0(n6525), .B1(
        image_data[487]), .Y(n6499) );
  AOI22XL U5319 ( .A0(n6524), .A1(image_data[295]), .B0(n6523), .B1(
        image_data[423]), .Y(n6500) );
  AOI22XL U5320 ( .A0(n6522), .A1(image_data[327]), .B0(n6521), .B1(
        image_data[455]), .Y(n6501) );
  AOI22XL U5321 ( .A0(n6520), .A1(image_data[263]), .B0(n6519), .B1(
        image_data[391]), .Y(n6502) );
  NAND4XL U5322 ( .A(n6554), .B(n6553), .C(n6552), .D(n6551), .Y(n6568) );
  AOI22XL U5323 ( .A0(n6544), .A1(image_data[15]), .B0(n6543), .B1(
        image_data[143]), .Y(n6554) );
  AOI22XL U5324 ( .A0(n6546), .A1(image_data[79]), .B0(n6545), .B1(
        image_data[207]), .Y(n6553) );
  AOI22XL U5325 ( .A0(n6548), .A1(image_data[47]), .B0(n6547), .B1(
        image_data[175]), .Y(n6552) );
  NAND4XL U5326 ( .A(n6566), .B(n6565), .C(n6564), .D(n6563), .Y(n6567) );
  AOI22XL U5327 ( .A0(n6556), .A1(image_data[31]), .B0(n6555), .B1(
        image_data[159]), .Y(n6566) );
  AOI22XL U5328 ( .A0(n6558), .A1(image_data[95]), .B0(n6557), .B1(
        image_data[223]), .Y(n6565) );
  AOI22XL U5329 ( .A0(n6560), .A1(image_data[63]), .B0(n6559), .B1(
        image_data[191]), .Y(n6564) );
  NAND4XL U5330 ( .A(n6542), .B(n6541), .C(n6540), .D(n6539), .Y(n6569) );
  AOI22XL U5331 ( .A0(n6532), .A1(image_data[23]), .B0(n6531), .B1(
        image_data[151]), .Y(n6542) );
  AOI22XL U5332 ( .A0(n6534), .A1(image_data[87]), .B0(n6533), .B1(
        image_data[215]), .Y(n6541) );
  AOI22XL U5333 ( .A0(n6536), .A1(image_data[55]), .B0(n6535), .B1(
        image_data[183]), .Y(n6540) );
  NAND4XL U5334 ( .A(n6530), .B(n6529), .C(n6528), .D(n6527), .Y(n6570) );
  AOI22XL U5335 ( .A0(n6520), .A1(image_data[7]), .B0(n6519), .B1(
        image_data[135]), .Y(n6530) );
  AOI22XL U5336 ( .A0(n6522), .A1(image_data[71]), .B0(n6521), .B1(
        image_data[199]), .Y(n6529) );
  AOI22XL U5337 ( .A0(n6524), .A1(image_data[39]), .B0(n6523), .B1(
        image_data[167]), .Y(n6528) );
  NAND4XL U5338 ( .A(n6510), .B(n6509), .C(n6508), .D(n6507), .Y(n6516) );
  AOI22XL U5339 ( .A0(n6544), .A1(image_data[271]), .B0(n6543), .B1(
        image_data[399]), .Y(n6510) );
  AOI22XL U5340 ( .A0(n6546), .A1(image_data[335]), .B0(n6545), .B1(
        image_data[463]), .Y(n6509) );
  AOI22XL U5341 ( .A0(n6548), .A1(image_data[303]), .B0(n6547), .B1(
        image_data[431]), .Y(n6508) );
  NAND4XL U5342 ( .A(n6514), .B(n6513), .C(n6512), .D(n6511), .Y(n6515) );
  AOI22XL U5343 ( .A0(n6556), .A1(image_data[287]), .B0(n6555), .B1(
        image_data[415]), .Y(n6514) );
  AOI22XL U5344 ( .A0(n6558), .A1(image_data[351]), .B0(n6557), .B1(
        image_data[479]), .Y(n6513) );
  AOI22XL U5345 ( .A0(n6560), .A1(image_data[319]), .B0(n6559), .B1(
        image_data[447]), .Y(n6512) );
  NAND4XL U5346 ( .A(n6506), .B(n6505), .C(n6504), .D(n6503), .Y(n6517) );
  AOI22XL U5347 ( .A0(n6532), .A1(image_data[279]), .B0(n6531), .B1(
        image_data[407]), .Y(n6506) );
  AOI22XL U5348 ( .A0(n6534), .A1(image_data[343]), .B0(n6533), .B1(
        image_data[471]), .Y(n6505) );
  AOI22XL U5349 ( .A0(n6536), .A1(image_data[311]), .B0(n6535), .B1(
        image_data[439]), .Y(n6504) );
  AOI22XL U5350 ( .A0(n6486), .A1(image_data[383]), .B0(n6485), .B1(
        image_data[511]), .Y(n6435) );
  AOI22XL U5351 ( .A0(n6484), .A1(image_data[319]), .B0(n6483), .B1(
        image_data[447]), .Y(n6436) );
  AOI22XL U5352 ( .A0(n6482), .A1(image_data[351]), .B0(n6481), .B1(
        image_data[479]), .Y(n6437) );
  AOI22XL U5353 ( .A0(n6480), .A1(image_data[287]), .B0(n6479), .B1(
        image_data[415]), .Y(n6438) );
  NAND4XL U5354 ( .A(n6478), .B(n6477), .C(n6476), .D(n6475), .Y(n6492) );
  AOI22XL U5355 ( .A0(n6468), .A1(image_data[15]), .B0(n6467), .B1(
        image_data[143]), .Y(n6478) );
  AOI22XL U5356 ( .A0(n6470), .A1(image_data[79]), .B0(n6469), .B1(
        image_data[207]), .Y(n6477) );
  AOI22XL U5357 ( .A0(n6472), .A1(image_data[47]), .B0(n6471), .B1(
        image_data[175]), .Y(n6476) );
  NAND4XL U5358 ( .A(n6466), .B(n6465), .C(n6464), .D(n6463), .Y(n6493) );
  AOI22XL U5359 ( .A0(n6456), .A1(image_data[23]), .B0(n6455), .B1(
        image_data[151]), .Y(n6466) );
  AOI22XL U5360 ( .A0(n6458), .A1(image_data[87]), .B0(n6457), .B1(
        image_data[215]), .Y(n6465) );
  AOI22XL U5361 ( .A0(n6460), .A1(image_data[55]), .B0(n6459), .B1(
        image_data[183]), .Y(n6464) );
  NAND4XL U5362 ( .A(n6454), .B(n6453), .C(n6452), .D(n6451), .Y(n6494) );
  AOI22XL U5363 ( .A0(n6444), .A1(image_data[7]), .B0(n6443), .B1(
        image_data[135]), .Y(n6454) );
  AOI22XL U5364 ( .A0(n6446), .A1(image_data[71]), .B0(n6445), .B1(
        image_data[199]), .Y(n6453) );
  AOI22XL U5365 ( .A0(n6448), .A1(image_data[39]), .B0(n6447), .B1(
        image_data[167]), .Y(n6452) );
  NAND4XL U5366 ( .A(n6490), .B(n6489), .C(n6488), .D(n6487), .Y(n6491) );
  AOI22XL U5367 ( .A0(n6480), .A1(image_data[31]), .B0(n6479), .B1(
        image_data[159]), .Y(n6490) );
  AOI22XL U5368 ( .A0(n6482), .A1(image_data[95]), .B0(n6481), .B1(
        image_data[223]), .Y(n6489) );
  AOI22XL U5369 ( .A0(n6484), .A1(image_data[63]), .B0(n6483), .B1(
        image_data[191]), .Y(n6488) );
  NAND4XL U5370 ( .A(n6434), .B(n6433), .C(n6432), .D(n6431), .Y(n6440) );
  AOI22XL U5371 ( .A0(n6468), .A1(image_data[271]), .B0(n6467), .B1(
        image_data[399]), .Y(n6434) );
  AOI22XL U5372 ( .A0(n6470), .A1(image_data[335]), .B0(n6469), .B1(
        image_data[463]), .Y(n6433) );
  AOI22XL U5373 ( .A0(n6472), .A1(image_data[303]), .B0(n6471), .B1(
        image_data[431]), .Y(n6432) );
  NAND4XL U5374 ( .A(n6430), .B(n6429), .C(n6428), .D(n6427), .Y(n6441) );
  AOI22XL U5375 ( .A0(n6456), .A1(image_data[279]), .B0(n6455), .B1(
        image_data[407]), .Y(n6430) );
  AOI22XL U5376 ( .A0(n6458), .A1(image_data[343]), .B0(n6457), .B1(
        image_data[471]), .Y(n6429) );
  AOI22XL U5377 ( .A0(n6460), .A1(image_data[311]), .B0(n6459), .B1(
        image_data[439]), .Y(n6428) );
  NAND4XL U5378 ( .A(n6426), .B(n6425), .C(n6424), .D(n6423), .Y(n6442) );
  AOI22XL U5379 ( .A0(n6444), .A1(image_data[263]), .B0(n6443), .B1(
        image_data[391]), .Y(n6426) );
  AOI22XL U5380 ( .A0(n6446), .A1(image_data[327]), .B0(n6445), .B1(
        image_data[455]), .Y(n6425) );
  AOI22XL U5381 ( .A0(n6448), .A1(image_data[295]), .B0(n6447), .B1(
        image_data[423]), .Y(n6424) );
  NAND4XL U5382 ( .A(n5721), .B(n5720), .C(n5719), .D(n5718), .Y(n5727) );
  AOI22XL U5383 ( .A0(n6468), .A1(image_data[268]), .B0(n6467), .B1(
        image_data[396]), .Y(n5721) );
  AOI22XL U5384 ( .A0(n6470), .A1(image_data[332]), .B0(n6469), .B1(
        image_data[460]), .Y(n5720) );
  AOI22XL U5385 ( .A0(n6472), .A1(image_data[300]), .B0(n6471), .B1(
        image_data[428]), .Y(n5719) );
  NAND4XL U5386 ( .A(n5717), .B(n5716), .C(n5715), .D(n5714), .Y(n5728) );
  AOI22XL U5387 ( .A0(n6456), .A1(image_data[276]), .B0(n6455), .B1(
        image_data[404]), .Y(n5717) );
  AOI22XL U5388 ( .A0(n6458), .A1(image_data[340]), .B0(n6457), .B1(
        image_data[468]), .Y(n5716) );
  AOI22XL U5389 ( .A0(n6460), .A1(image_data[308]), .B0(n6459), .B1(
        image_data[436]), .Y(n5715) );
  NAND4XL U5390 ( .A(n5713), .B(n5712), .C(n5711), .D(n5710), .Y(n5729) );
  AOI22XL U5391 ( .A0(n6444), .A1(image_data[260]), .B0(n6443), .B1(
        image_data[388]), .Y(n5713) );
  AOI22XL U5392 ( .A0(n6446), .A1(image_data[324]), .B0(n6445), .B1(
        image_data[452]), .Y(n5712) );
  AOI22XL U5393 ( .A0(n6448), .A1(image_data[292]), .B0(n6447), .B1(
        image_data[420]), .Y(n5711) );
  NAND4XL U5394 ( .A(n5725), .B(n5724), .C(n5723), .D(n5722), .Y(n5726) );
  AOI22XL U5395 ( .A0(n6480), .A1(image_data[284]), .B0(n6479), .B1(
        image_data[412]), .Y(n5725) );
  AOI22XL U5396 ( .A0(n6482), .A1(image_data[348]), .B0(n6481), .B1(
        image_data[476]), .Y(n5724) );
  AOI22XL U5397 ( .A0(n6484), .A1(image_data[316]), .B0(n6483), .B1(
        image_data[444]), .Y(n5723) );
  NOR4XL U5398 ( .A(n5791), .B(n5790), .C(n5789), .D(n5788), .Y(n5792) );
  NAND4XL U5399 ( .A(n5787), .B(n5786), .C(n5785), .D(n5784), .Y(n5788) );
  NAND4XL U5400 ( .A(n5775), .B(n5774), .C(n5773), .D(n5772), .Y(n5791) );
  NAND4XL U5401 ( .A(n5779), .B(n5778), .C(n5777), .D(n5776), .Y(n5790) );
  NOR4XL U5402 ( .A(n5771), .B(n5770), .C(n5769), .D(n5768), .Y(n5793) );
  NAND4XL U5403 ( .A(n5767), .B(n5766), .C(n5765), .D(n5764), .Y(n5768) );
  NAND4XL U5404 ( .A(n5755), .B(n5754), .C(n5753), .D(n5752), .Y(n5771) );
  NAND4XL U5405 ( .A(n5759), .B(n5758), .C(n5757), .D(n5756), .Y(n5770) );
  NOR4XL U5406 ( .A(n5749), .B(n5748), .C(n5747), .D(n5746), .Y(n5750) );
  NAND4XL U5407 ( .A(n5745), .B(n5744), .C(n5743), .D(n5742), .Y(n5746) );
  NAND4XL U5408 ( .A(n5733), .B(n5732), .C(n5731), .D(n5730), .Y(n5749) );
  NAND4XL U5409 ( .A(n5737), .B(n5736), .C(n5735), .D(n5734), .Y(n5748) );
  AOI22XL U5410 ( .A0(n6486), .A1(image_data[122]), .B0(n6485), .B1(
        image_data[250]), .Y(n5073) );
  AOI22XL U5411 ( .A0(n6484), .A1(image_data[58]), .B0(n6483), .B1(
        image_data[186]), .Y(n5074) );
  AOI22XL U5412 ( .A0(n6482), .A1(image_data[90]), .B0(n6481), .B1(
        image_data[218]), .Y(n5075) );
  AOI22XL U5413 ( .A0(n6480), .A1(image_data[26]), .B0(n6479), .B1(
        image_data[154]), .Y(n5076) );
  AOI22XL U5414 ( .A0(n6450), .A1(image_data[98]), .B0(n6449), .B1(
        image_data[226]), .Y(n5061) );
  AOI22XL U5415 ( .A0(n6448), .A1(image_data[34]), .B0(n6447), .B1(
        image_data[162]), .Y(n5062) );
  AOI22XL U5416 ( .A0(n6446), .A1(image_data[66]), .B0(n6445), .B1(
        image_data[194]), .Y(n5063) );
  AOI22XL U5417 ( .A0(n6444), .A1(image_data[2]), .B0(n6443), .B1(
        image_data[130]), .Y(n5064) );
  AOI22XL U5418 ( .A0(n6462), .A1(image_data[114]), .B0(n6461), .B1(
        image_data[242]), .Y(n5065) );
  AOI22XL U5419 ( .A0(n6460), .A1(image_data[50]), .B0(n6459), .B1(
        image_data[178]), .Y(n5066) );
  AOI22XL U5420 ( .A0(n6458), .A1(image_data[82]), .B0(n6457), .B1(
        image_data[210]), .Y(n5067) );
  AOI22XL U5421 ( .A0(n6456), .A1(image_data[18]), .B0(n6455), .B1(
        image_data[146]), .Y(n5068) );
  NAND4XL U5422 ( .A(n5072), .B(n5071), .C(n5070), .D(n5069), .Y(n5078) );
  AOI22XL U5423 ( .A0(n6468), .A1(image_data[10]), .B0(n6467), .B1(
        image_data[138]), .Y(n5072) );
  AOI22XL U5424 ( .A0(n6470), .A1(image_data[74]), .B0(n6469), .B1(
        image_data[202]), .Y(n5071) );
  AOI22XL U5425 ( .A0(n6472), .A1(image_data[42]), .B0(n6471), .B1(
        image_data[170]), .Y(n5070) );
  AOI22XL U5426 ( .A0(n6486), .A1(image_data[378]), .B0(n6485), .B1(
        image_data[506]), .Y(n5053) );
  AOI22XL U5427 ( .A0(n6484), .A1(image_data[314]), .B0(n6483), .B1(
        image_data[442]), .Y(n5054) );
  AOI22XL U5428 ( .A0(n6482), .A1(image_data[346]), .B0(n6481), .B1(
        image_data[474]), .Y(n5055) );
  AOI22XL U5429 ( .A0(n6480), .A1(image_data[282]), .B0(n6479), .B1(
        image_data[410]), .Y(n5056) );
  AOI22XL U5430 ( .A0(n6450), .A1(image_data[354]), .B0(n6449), .B1(
        image_data[482]), .Y(n5026) );
  AOI22XL U5431 ( .A0(n6448), .A1(image_data[290]), .B0(n6447), .B1(
        image_data[418]), .Y(n5027) );
  AOI22XL U5432 ( .A0(n6446), .A1(image_data[322]), .B0(n6445), .B1(
        image_data[450]), .Y(n5028) );
  AOI22XL U5433 ( .A0(n6444), .A1(image_data[258]), .B0(n6443), .B1(
        image_data[386]), .Y(n5029) );
  AOI22XL U5434 ( .A0(n6462), .A1(image_data[370]), .B0(n6461), .B1(
        image_data[498]), .Y(n5032) );
  AOI22XL U5435 ( .A0(n6460), .A1(image_data[306]), .B0(n6459), .B1(
        image_data[434]), .Y(n5033) );
  AOI22XL U5436 ( .A0(n6458), .A1(image_data[338]), .B0(n6457), .B1(
        image_data[466]), .Y(n5034) );
  AOI22XL U5437 ( .A0(n6456), .A1(image_data[274]), .B0(n6455), .B1(
        image_data[402]), .Y(n5035) );
  NAND4XL U5438 ( .A(n5041), .B(n5040), .C(n5039), .D(n5038), .Y(n5058) );
  AOI22XL U5439 ( .A0(n6468), .A1(image_data[266]), .B0(n6467), .B1(
        image_data[394]), .Y(n5041) );
  AOI22XL U5440 ( .A0(n6470), .A1(image_data[330]), .B0(n6469), .B1(
        image_data[458]), .Y(n5040) );
  AOI22XL U5441 ( .A0(n6472), .A1(image_data[298]), .B0(n6471), .B1(
        image_data[426]), .Y(n5039) );
  AOI22XL U5442 ( .A0(n6534), .A1(image_data[338]), .B0(n6533), .B1(
        image_data[466]), .Y(n5206) );
  AOI22XL U5443 ( .A0(n6538), .A1(image_data[370]), .B0(n6537), .B1(
        image_data[498]), .Y(n5204) );
  AOI22XL U5444 ( .A0(n6536), .A1(image_data[306]), .B0(n6535), .B1(
        image_data[434]), .Y(n5205) );
  AOI22XL U5445 ( .A0(n6532), .A1(image_data[274]), .B0(n6531), .B1(
        image_data[402]), .Y(n5207) );
  NAND4XL U5446 ( .A(n5244), .B(n5243), .C(n5242), .D(n5241), .Y(n5250) );
  AOI22XL U5447 ( .A0(n6544), .A1(image_data[10]), .B0(n6543), .B1(
        image_data[138]), .Y(n5244) );
  AOI22XL U5448 ( .A0(n6546), .A1(image_data[74]), .B0(n6545), .B1(
        image_data[202]), .Y(n5243) );
  AOI22XL U5449 ( .A0(n6548), .A1(image_data[42]), .B0(n6547), .B1(
        image_data[170]), .Y(n5242) );
  NAND4XL U5450 ( .A(n5248), .B(n5247), .C(n5246), .D(n5245), .Y(n5249) );
  AOI22XL U5451 ( .A0(n6556), .A1(image_data[26]), .B0(n6555), .B1(
        image_data[154]), .Y(n5248) );
  AOI22XL U5452 ( .A0(n6558), .A1(image_data[90]), .B0(n6557), .B1(
        image_data[218]), .Y(n5247) );
  AOI22XL U5453 ( .A0(n6560), .A1(image_data[58]), .B0(n6559), .B1(
        image_data[186]), .Y(n5246) );
  NAND4XL U5454 ( .A(n5236), .B(n5235), .C(n5234), .D(n5233), .Y(n5252) );
  AOI22XL U5455 ( .A0(n6520), .A1(image_data[2]), .B0(n6519), .B1(
        image_data[130]), .Y(n5236) );
  AOI22XL U5456 ( .A0(n6522), .A1(image_data[66]), .B0(n6521), .B1(
        image_data[194]), .Y(n5235) );
  AOI22XL U5457 ( .A0(n6524), .A1(image_data[34]), .B0(n6523), .B1(
        image_data[162]), .Y(n5234) );
  NAND4XL U5458 ( .A(n5240), .B(n5239), .C(n5238), .D(n5237), .Y(n5251) );
  AOI22XL U5459 ( .A0(n6532), .A1(image_data[18]), .B0(n6531), .B1(
        image_data[146]), .Y(n5240) );
  AOI22XL U5460 ( .A0(n6536), .A1(image_data[50]), .B0(n6535), .B1(
        image_data[178]), .Y(n5238) );
  AOI22XL U5461 ( .A0(n6538), .A1(image_data[114]), .B0(n6537), .B1(
        image_data[242]), .Y(n5237) );
  NAND4XL U5462 ( .A(n5213), .B(n5212), .C(n5211), .D(n5210), .Y(n5230) );
  AOI22XL U5463 ( .A0(n6544), .A1(image_data[266]), .B0(n6543), .B1(
        image_data[394]), .Y(n5213) );
  AOI22XL U5464 ( .A0(n6546), .A1(image_data[330]), .B0(n6545), .B1(
        image_data[458]), .Y(n5212) );
  AOI22XL U5465 ( .A0(n6548), .A1(image_data[298]), .B0(n6547), .B1(
        image_data[426]), .Y(n5211) );
  NAND4XL U5466 ( .A(n5228), .B(n5227), .C(n5226), .D(n5225), .Y(n5229) );
  AOI22XL U5467 ( .A0(n6556), .A1(image_data[282]), .B0(n6555), .B1(
        image_data[410]), .Y(n5228) );
  AOI22XL U5468 ( .A0(n6558), .A1(image_data[346]), .B0(n6557), .B1(
        image_data[474]), .Y(n5227) );
  AOI22XL U5469 ( .A0(n6560), .A1(image_data[314]), .B0(n6559), .B1(
        image_data[442]), .Y(n5226) );
  NAND4XL U5470 ( .A(n5201), .B(n5200), .C(n5199), .D(n5198), .Y(n5232) );
  AOI22XL U5471 ( .A0(n6520), .A1(image_data[258]), .B0(n6519), .B1(
        image_data[386]), .Y(n5201) );
  AOI22XL U5472 ( .A0(n6522), .A1(image_data[322]), .B0(n6521), .B1(
        image_data[450]), .Y(n5200) );
  AOI22XL U5473 ( .A0(n6524), .A1(image_data[290]), .B0(n6523), .B1(
        image_data[418]), .Y(n5199) );
  AOI22X1 U5474 ( .A0(n3450), .A1(n3821), .B0(n3820), .B1(n4959), .Y(N2760) );
  NOR4XL U5475 ( .A(n3790), .B(n3789), .C(n3788), .D(n3787), .Y(n3821) );
  NOR4XL U5476 ( .A(n3819), .B(n3818), .C(n3817), .D(n3816), .Y(n3820) );
  NAND4XL U5477 ( .A(n3778), .B(n3777), .C(n3776), .D(n3775), .Y(n3789) );
  AOI22XL U5478 ( .A0(n3935), .A1(image_data[373]), .B0(n3888), .B1(
        image_data[501]), .Y(n4497) );
  AOI22XL U5479 ( .A0(n3887), .A1(image_data[309]), .B0(n3936), .B1(
        image_data[437]), .Y(n4498) );
  AOI22XL U5480 ( .A0(n3884), .A1(image_data[277]), .B0(n3934), .B1(
        image_data[405]), .Y(n4500) );
  AOI22XL U5481 ( .A0(n3885), .A1(image_data[341]), .B0(n3886), .B1(
        image_data[469]), .Y(n4499) );
  NAND4XL U5482 ( .A(n4516), .B(n4515), .C(n4514), .D(n4513), .Y(n4532) );
  AOI22XL U5483 ( .A0(n3897), .A1(image_data[5]), .B0(n3896), .B1(
        image_data[133]), .Y(n4516) );
  AOI22XL U5484 ( .A0(n3928), .A1(image_data[37]), .B0(n3929), .B1(
        image_data[165]), .Y(n4514) );
  AOI22XL U5485 ( .A0(n3893), .A1(image_data[101]), .B0(n3894), .B1(
        image_data[229]), .Y(n4513) );
  NAND4XL U5486 ( .A(n4528), .B(n4527), .C(n4526), .D(n4525), .Y(n4529) );
  AOI22XL U5487 ( .A0(n3875), .A1(image_data[93]), .B0(n3876), .B1(
        image_data[221]), .Y(n4527) );
  AOI22XL U5488 ( .A0(n3877), .A1(image_data[61]), .B0(n3949), .B1(
        image_data[189]), .Y(n4526) );
  AOI22XL U5489 ( .A0(n3874), .A1(image_data[29]), .B0(n3948), .B1(
        image_data[157]), .Y(n4528) );
  NAND4XL U5490 ( .A(n4524), .B(n4523), .C(n4522), .D(n4521), .Y(n4530) );
  AOI22XL U5491 ( .A0(n3866), .A1(image_data[77]), .B0(n3867), .B1(
        image_data[205]), .Y(n4523) );
  AOI22XL U5492 ( .A0(n3865), .A1(image_data[13]), .B0(n3941), .B1(
        image_data[141]), .Y(n4524) );
  AOI22XL U5493 ( .A0(n3942), .A1(image_data[45]), .B0(n3943), .B1(
        image_data[173]), .Y(n4522) );
  NAND4XL U5494 ( .A(n4520), .B(n4519), .C(n4518), .D(n4517), .Y(n4531) );
  AOI22XL U5495 ( .A0(n3885), .A1(image_data[85]), .B0(n3886), .B1(
        image_data[213]), .Y(n4519) );
  AOI22XL U5496 ( .A0(n3884), .A1(image_data[21]), .B0(n3934), .B1(
        image_data[149]), .Y(n4520) );
  AOI22XL U5497 ( .A0(n3887), .A1(image_data[53]), .B0(n3936), .B1(
        image_data[181]), .Y(n4518) );
  NAND4XL U5498 ( .A(n4496), .B(n4495), .C(n4494), .D(n4493), .Y(n4512) );
  AOI22XL U5499 ( .A0(n3897), .A1(image_data[261]), .B0(n3896), .B1(
        image_data[389]), .Y(n4496) );
  AOI22XL U5500 ( .A0(n3928), .A1(image_data[293]), .B0(n3929), .B1(
        image_data[421]), .Y(n4494) );
  AOI22XL U5501 ( .A0(n3893), .A1(image_data[357]), .B0(n3894), .B1(
        image_data[485]), .Y(n4493) );
  NAND4XL U5502 ( .A(n4508), .B(n4507), .C(n4506), .D(n4505), .Y(n4509) );
  AOI22XL U5503 ( .A0(n3875), .A1(image_data[349]), .B0(n3876), .B1(
        image_data[477]), .Y(n4507) );
  AOI22XL U5504 ( .A0(n3877), .A1(image_data[317]), .B0(n3949), .B1(
        image_data[445]), .Y(n4506) );
  AOI22XL U5505 ( .A0(n3874), .A1(image_data[285]), .B0(n3948), .B1(
        image_data[413]), .Y(n4508) );
  NAND4XL U5506 ( .A(n4504), .B(n4503), .C(n4502), .D(n4501), .Y(n4510) );
  AOI22XL U5507 ( .A0(n3866), .A1(image_data[333]), .B0(n3867), .B1(
        image_data[461]), .Y(n4503) );
  AOI22XL U5508 ( .A0(n3865), .A1(image_data[269]), .B0(n3941), .B1(
        image_data[397]), .Y(n4504) );
  AOI22XL U5509 ( .A0(n3942), .A1(image_data[301]), .B0(n3943), .B1(
        image_data[429]), .Y(n4502) );
  AOI22XL U5510 ( .A0(n3869), .A1(image_data[293]), .B0(n3868), .B1(
        image_data[421]), .Y(n3519) );
  AOI22XL U5511 ( .A0(n3942), .A1(image_data[357]), .B0(n3943), .B1(
        image_data[485]), .Y(n3518) );
  AOI22XL U5512 ( .A0(n3865), .A1(image_data[325]), .B0(n3941), .B1(
        image_data[453]), .Y(n3520) );
  AOI22XL U5513 ( .A0(n3867), .A1(image_data[261]), .B0(n3866), .B1(
        image_data[389]), .Y(n3521) );
  NAND4XL U5514 ( .A(n3553), .B(n3552), .C(n3551), .D(n3550), .Y(n3554) );
  AOI22XL U5515 ( .A0(n3897), .A1(image_data[61]), .B0(n3896), .B1(
        image_data[189]), .Y(n3551) );
  AOI22XL U5516 ( .A0(n3928), .A1(image_data[93]), .B0(n3929), .B1(
        image_data[221]), .Y(n3552) );
  AOI22XL U5517 ( .A0(n3894), .A1(image_data[29]), .B0(n3893), .B1(
        image_data[157]), .Y(n3553) );
  NAND4XL U5518 ( .A(n3549), .B(n3548), .C(n3547), .D(n3546), .Y(n3555) );
  AOI22XL U5519 ( .A0(n3886), .A1(image_data[13]), .B0(n3885), .B1(
        image_data[141]), .Y(n3549) );
  AOI22XL U5520 ( .A0(n3887), .A1(image_data[109]), .B0(n3936), .B1(
        image_data[237]), .Y(n3546) );
  AOI22XL U5521 ( .A0(n3884), .A1(image_data[77]), .B0(n3934), .B1(
        image_data[205]), .Y(n3548) );
  NAND4XL U5522 ( .A(n3545), .B(n3544), .C(n3543), .D(n3542), .Y(n3556) );
  AOI22XL U5523 ( .A0(n3876), .A1(image_data[21]), .B0(n3875), .B1(
        image_data[149]), .Y(n3545) );
  AOI22XL U5524 ( .A0(n3877), .A1(image_data[117]), .B0(n3949), .B1(
        image_data[245]), .Y(n3542) );
  AOI22XL U5525 ( .A0(n3874), .A1(image_data[85]), .B0(n3948), .B1(
        image_data[213]), .Y(n3544) );
  NAND4XL U5526 ( .A(n3541), .B(n3540), .C(n3539), .D(n3538), .Y(n3557) );
  AOI22XL U5527 ( .A0(n3867), .A1(image_data[5]), .B0(n3866), .B1(
        image_data[133]), .Y(n3541) );
  AOI22XL U5528 ( .A0(n3865), .A1(image_data[69]), .B0(n3941), .B1(
        image_data[197]), .Y(n3540) );
  AOI22XL U5529 ( .A0(n3942), .A1(image_data[101]), .B0(n3943), .B1(
        image_data[229]), .Y(n3538) );
  NAND4XL U5530 ( .A(n3533), .B(n3532), .C(n3531), .D(n3530), .Y(n3534) );
  AOI22XL U5531 ( .A0(n3897), .A1(image_data[317]), .B0(n3896), .B1(
        image_data[445]), .Y(n3531) );
  AOI22XL U5532 ( .A0(n3928), .A1(image_data[349]), .B0(n3929), .B1(
        image_data[477]), .Y(n3532) );
  AOI22XL U5533 ( .A0(n3894), .A1(image_data[285]), .B0(n3893), .B1(
        image_data[413]), .Y(n3533) );
  NAND4XL U5534 ( .A(n3529), .B(n3528), .C(n3527), .D(n3526), .Y(n3535) );
  AOI22XL U5535 ( .A0(n3886), .A1(image_data[269]), .B0(n3885), .B1(
        image_data[397]), .Y(n3529) );
  AOI22XL U5536 ( .A0(n3887), .A1(image_data[365]), .B0(n3936), .B1(
        image_data[493]), .Y(n3526) );
  AOI22XL U5537 ( .A0(n3884), .A1(image_data[333]), .B0(n3934), .B1(
        image_data[461]), .Y(n3528) );
  NAND4XL U5538 ( .A(n3525), .B(n3524), .C(n3523), .D(n3522), .Y(n3536) );
  AOI22XL U5539 ( .A0(n3876), .A1(image_data[277]), .B0(n3875), .B1(
        image_data[405]), .Y(n3525) );
  AOI22XL U5540 ( .A0(n3877), .A1(image_data[373]), .B0(n3949), .B1(
        image_data[501]), .Y(n3522) );
  AOI22XL U5541 ( .A0(n3874), .A1(image_data[341]), .B0(n3948), .B1(
        image_data[469]), .Y(n3524) );
  AOI22XL U5542 ( .A0(n3884), .A1(image_data[276]), .B0(n3934), .B1(
        image_data[404]), .Y(n4458) );
  AOI22XL U5543 ( .A0(n3885), .A1(image_data[340]), .B0(n3886), .B1(
        image_data[468]), .Y(n4457) );
  NOR2XL U5544 ( .A(n5706), .B(n4588), .Y(n6281) );
  AOI22XL U5545 ( .A0(n6562), .A1(image_data[381]), .B0(n6561), .B1(
        image_data[509]), .Y(n5985) );
  AOI22XL U5546 ( .A0(n6560), .A1(image_data[317]), .B0(n6559), .B1(
        image_data[445]), .Y(n5986) );
  AOI22XL U5547 ( .A0(n6558), .A1(image_data[349]), .B0(n6557), .B1(
        image_data[477]), .Y(n5987) );
  AOI22XL U5548 ( .A0(n6556), .A1(image_data[285]), .B0(n6555), .B1(
        image_data[413]), .Y(n5988) );
  NAND4XL U5549 ( .A(n6004), .B(n6003), .C(n6002), .D(n6001), .Y(n6010) );
  AOI22XL U5550 ( .A0(n6544), .A1(image_data[13]), .B0(n6543), .B1(
        image_data[141]), .Y(n6004) );
  AOI22XL U5551 ( .A0(n6546), .A1(image_data[77]), .B0(n6545), .B1(
        image_data[205]), .Y(n6003) );
  AOI22XL U5552 ( .A0(n6548), .A1(image_data[45]), .B0(n6547), .B1(
        image_data[173]), .Y(n6002) );
  NAND4XL U5553 ( .A(n6000), .B(n5999), .C(n5998), .D(n5997), .Y(n6011) );
  AOI22XL U5554 ( .A0(n6532), .A1(image_data[21]), .B0(n6531), .B1(
        image_data[149]), .Y(n6000) );
  AOI22XL U5555 ( .A0(n6534), .A1(image_data[85]), .B0(n6533), .B1(
        image_data[213]), .Y(n5999) );
  AOI22XL U5556 ( .A0(n6536), .A1(image_data[53]), .B0(n6535), .B1(
        image_data[181]), .Y(n5998) );
  NAND4XL U5557 ( .A(n5996), .B(n5995), .C(n5994), .D(n5993), .Y(n6012) );
  AOI22XL U5558 ( .A0(n6520), .A1(image_data[5]), .B0(n6519), .B1(
        image_data[133]), .Y(n5996) );
  AOI22XL U5559 ( .A0(n6522), .A1(image_data[69]), .B0(n6521), .B1(
        image_data[197]), .Y(n5995) );
  AOI22XL U5560 ( .A0(n6524), .A1(image_data[37]), .B0(n6523), .B1(
        image_data[165]), .Y(n5994) );
  NAND4XL U5561 ( .A(n6008), .B(n6007), .C(n6006), .D(n6005), .Y(n6009) );
  AOI22XL U5562 ( .A0(n6556), .A1(image_data[29]), .B0(n6555), .B1(
        image_data[157]), .Y(n6008) );
  AOI22XL U5563 ( .A0(n6558), .A1(image_data[93]), .B0(n6557), .B1(
        image_data[221]), .Y(n6007) );
  AOI22XL U5564 ( .A0(n6560), .A1(image_data[61]), .B0(n6559), .B1(
        image_data[189]), .Y(n6006) );
  NAND4XL U5565 ( .A(n5984), .B(n5983), .C(n5982), .D(n5981), .Y(n5990) );
  AOI22XL U5566 ( .A0(n6544), .A1(image_data[269]), .B0(n6543), .B1(
        image_data[397]), .Y(n5984) );
  AOI22XL U5567 ( .A0(n6546), .A1(image_data[333]), .B0(n6545), .B1(
        image_data[461]), .Y(n5983) );
  AOI22XL U5568 ( .A0(n6548), .A1(image_data[301]), .B0(n6547), .B1(
        image_data[429]), .Y(n5982) );
  NAND4XL U5569 ( .A(n5980), .B(n5979), .C(n5978), .D(n5977), .Y(n5991) );
  AOI22XL U5570 ( .A0(n6532), .A1(image_data[277]), .B0(n6531), .B1(
        image_data[405]), .Y(n5980) );
  AOI22XL U5571 ( .A0(n6534), .A1(image_data[341]), .B0(n6533), .B1(
        image_data[469]), .Y(n5979) );
  AOI22XL U5572 ( .A0(n6536), .A1(image_data[309]), .B0(n6535), .B1(
        image_data[437]), .Y(n5978) );
  NAND4XL U5573 ( .A(n5976), .B(n5975), .C(n5974), .D(n5973), .Y(n5992) );
  AOI22XL U5574 ( .A0(n6520), .A1(image_data[261]), .B0(n6519), .B1(
        image_data[389]), .Y(n5976) );
  AOI22XL U5575 ( .A0(n6522), .A1(image_data[325]), .B0(n6521), .B1(
        image_data[453]), .Y(n5975) );
  AOI22XL U5576 ( .A0(n6524), .A1(image_data[293]), .B0(n6523), .B1(
        image_data[421]), .Y(n5974) );
  AOI22XL U5577 ( .A0(n3465), .A1(n5185), .B0(n5187), .B1(n3450), .Y(n5169) );
  AOI22XL U5578 ( .A0(op4[5]), .A1(n5183), .B0(n5182), .B1(n5165), .Y(n5170)
         );
  AOI22XL U5579 ( .A0(n6486), .A1(image_data[381]), .B0(n6485), .B1(
        image_data[509]), .Y(n5943) );
  AOI22XL U5580 ( .A0(n6484), .A1(image_data[317]), .B0(n6483), .B1(
        image_data[445]), .Y(n5944) );
  AOI22XL U5581 ( .A0(n6482), .A1(image_data[349]), .B0(n6481), .B1(
        image_data[477]), .Y(n5945) );
  AOI22XL U5582 ( .A0(n6480), .A1(image_data[285]), .B0(n6479), .B1(
        image_data[413]), .Y(n5946) );
  NAND4XL U5583 ( .A(n5962), .B(n5961), .C(n5960), .D(n5959), .Y(n5968) );
  AOI22XL U5584 ( .A0(n6468), .A1(image_data[13]), .B0(n6467), .B1(
        image_data[141]), .Y(n5962) );
  AOI22XL U5585 ( .A0(n6470), .A1(image_data[77]), .B0(n6469), .B1(
        image_data[205]), .Y(n5961) );
  AOI22XL U5586 ( .A0(n6472), .A1(image_data[45]), .B0(n6471), .B1(
        image_data[173]), .Y(n5960) );
  NAND4XL U5587 ( .A(n5958), .B(n5957), .C(n5956), .D(n5955), .Y(n5969) );
  AOI22XL U5588 ( .A0(n6456), .A1(image_data[21]), .B0(n6455), .B1(
        image_data[149]), .Y(n5958) );
  AOI22XL U5589 ( .A0(n6458), .A1(image_data[85]), .B0(n6457), .B1(
        image_data[213]), .Y(n5957) );
  AOI22XL U5590 ( .A0(n6460), .A1(image_data[53]), .B0(n6459), .B1(
        image_data[181]), .Y(n5956) );
  NAND4XL U5591 ( .A(n5954), .B(n5953), .C(n5952), .D(n5951), .Y(n5970) );
  AOI22XL U5592 ( .A0(n6444), .A1(image_data[5]), .B0(n6443), .B1(
        image_data[133]), .Y(n5954) );
  AOI22XL U5593 ( .A0(n6446), .A1(image_data[69]), .B0(n6445), .B1(
        image_data[197]), .Y(n5953) );
  AOI22XL U5594 ( .A0(n6448), .A1(image_data[37]), .B0(n6447), .B1(
        image_data[165]), .Y(n5952) );
  NAND4XL U5595 ( .A(n5966), .B(n5965), .C(n5964), .D(n5963), .Y(n5967) );
  AOI22XL U5596 ( .A0(n6480), .A1(image_data[29]), .B0(n6479), .B1(
        image_data[157]), .Y(n5966) );
  AOI22XL U5597 ( .A0(n6482), .A1(image_data[93]), .B0(n6481), .B1(
        image_data[221]), .Y(n5965) );
  AOI22XL U5598 ( .A0(n6484), .A1(image_data[61]), .B0(n6483), .B1(
        image_data[189]), .Y(n5964) );
  NAND4XL U5599 ( .A(n5942), .B(n5941), .C(n5940), .D(n5939), .Y(n5948) );
  AOI22XL U5600 ( .A0(n6468), .A1(image_data[269]), .B0(n6467), .B1(
        image_data[397]), .Y(n5942) );
  AOI22XL U5601 ( .A0(n6470), .A1(image_data[333]), .B0(n6469), .B1(
        image_data[461]), .Y(n5941) );
  AOI22XL U5602 ( .A0(n6472), .A1(image_data[301]), .B0(n6471), .B1(
        image_data[429]), .Y(n5940) );
  NAND4XL U5603 ( .A(n5938), .B(n5937), .C(n5936), .D(n5935), .Y(n5949) );
  AOI22XL U5604 ( .A0(n6456), .A1(image_data[277]), .B0(n6455), .B1(
        image_data[405]), .Y(n5938) );
  AOI22XL U5605 ( .A0(n6458), .A1(image_data[341]), .B0(n6457), .B1(
        image_data[469]), .Y(n5937) );
  AOI22XL U5606 ( .A0(n6460), .A1(image_data[309]), .B0(n6459), .B1(
        image_data[437]), .Y(n5936) );
  NAND4XL U5607 ( .A(n5934), .B(n5933), .C(n5932), .D(n5931), .Y(n5950) );
  AOI22XL U5608 ( .A0(n6444), .A1(image_data[261]), .B0(n6443), .B1(
        image_data[389]), .Y(n5934) );
  AOI22XL U5609 ( .A0(n6446), .A1(image_data[325]), .B0(n6445), .B1(
        image_data[453]), .Y(n5933) );
  AOI22XL U5610 ( .A0(n6448), .A1(image_data[293]), .B0(n6447), .B1(
        image_data[421]), .Y(n5932) );
  CMPR32X1 U5611 ( .A(DP_OP_2677J1_122_9848_n15), .B(DP_OP_2677J1_122_9848_n17), .C(n5897), .CO(n6015), .S(n5795) );
  AOI22XL U5612 ( .A0(n3935), .A1(image_data[374]), .B0(n3888), .B1(
        image_data[502]), .Y(n4406) );
  AOI22XL U5613 ( .A0(n3884), .A1(image_data[278]), .B0(n4427), .B1(
        image_data[406]), .Y(n4409) );
  AOI22XL U5614 ( .A0(n3887), .A1(image_data[310]), .B0(n4428), .B1(
        image_data[438]), .Y(n4407) );
  AOI22XL U5615 ( .A0(n3885), .A1(image_data[342]), .B0(n3886), .B1(
        image_data[470]), .Y(n4408) );
  NAND4XL U5616 ( .A(n4426), .B(n4425), .C(n4424), .D(n4423), .Y(n4448) );
  AOI22XL U5617 ( .A0(n3897), .A1(image_data[6]), .B0(n3896), .B1(
        image_data[134]), .Y(n4426) );
  AOI22XL U5618 ( .A0(n3928), .A1(image_data[38]), .B0(n4422), .B1(
        image_data[166]), .Y(n4424) );
  AOI22XL U5619 ( .A0(n3893), .A1(image_data[102]), .B0(n3894), .B1(
        image_data[230]), .Y(n4423) );
  NAND4XL U5620 ( .A(n4444), .B(n4443), .C(n4442), .D(n4441), .Y(n4445) );
  AOI22XL U5621 ( .A0(n3875), .A1(image_data[94]), .B0(n3876), .B1(
        image_data[222]), .Y(n4443) );
  AOI22XL U5622 ( .A0(n3874), .A1(image_data[30]), .B0(n4439), .B1(
        image_data[158]), .Y(n4444) );
  AOI22XL U5623 ( .A0(n3877), .A1(image_data[62]), .B0(n4440), .B1(
        image_data[190]), .Y(n4442) );
  NAND4XL U5624 ( .A(n4438), .B(n4437), .C(n4436), .D(n4435), .Y(n4446) );
  AOI22XL U5625 ( .A0(n3865), .A1(image_data[14]), .B0(n4433), .B1(
        image_data[142]), .Y(n4438) );
  AOI22XL U5626 ( .A0(n3866), .A1(image_data[78]), .B0(n3867), .B1(
        image_data[206]), .Y(n4437) );
  AOI22XL U5627 ( .A0(n3942), .A1(image_data[46]), .B0(n4434), .B1(
        image_data[174]), .Y(n4436) );
  NAND4XL U5628 ( .A(n4432), .B(n4431), .C(n4430), .D(n4429), .Y(n4447) );
  AOI22XL U5629 ( .A0(n3885), .A1(image_data[86]), .B0(n3886), .B1(
        image_data[214]), .Y(n4431) );
  AOI22XL U5630 ( .A0(n3887), .A1(image_data[54]), .B0(n4428), .B1(
        image_data[182]), .Y(n4430) );
  AOI22XL U5631 ( .A0(n3884), .A1(image_data[22]), .B0(n4427), .B1(
        image_data[150]), .Y(n4432) );
  NAND4XL U5632 ( .A(n4405), .B(n4404), .C(n4403), .D(n4402), .Y(n4421) );
  AOI22XL U5633 ( .A0(n3928), .A1(image_data[294]), .B0(n4422), .B1(
        image_data[422]), .Y(n4403) );
  AOI22XL U5634 ( .A0(n3897), .A1(image_data[262]), .B0(n3896), .B1(
        image_data[390]), .Y(n4405) );
  AOI22XL U5635 ( .A0(n3893), .A1(image_data[358]), .B0(n3894), .B1(
        image_data[486]), .Y(n4402) );
  NAND4XL U5636 ( .A(n4417), .B(n4416), .C(n4415), .D(n4414), .Y(n4418) );
  AOI22XL U5637 ( .A0(n3875), .A1(image_data[350]), .B0(n3876), .B1(
        image_data[478]), .Y(n4416) );
  AOI22XL U5638 ( .A0(n3874), .A1(image_data[286]), .B0(n4439), .B1(
        image_data[414]), .Y(n4417) );
  AOI22XL U5639 ( .A0(n3877), .A1(image_data[318]), .B0(n4440), .B1(
        image_data[446]), .Y(n4415) );
  NAND4XL U5640 ( .A(n4413), .B(n4412), .C(n4411), .D(n4410), .Y(n4419) );
  AOI22XL U5641 ( .A0(n3866), .A1(image_data[334]), .B0(n3867), .B1(
        image_data[462]), .Y(n4412) );
  AOI22XL U5642 ( .A0(n3865), .A1(image_data[270]), .B0(n4433), .B1(
        image_data[398]), .Y(n4413) );
  AOI22XL U5643 ( .A0(n3942), .A1(image_data[302]), .B0(n4434), .B1(
        image_data[430]), .Y(n4411) );
  AOI22XL U5644 ( .A0(n3869), .A1(image_data[294]), .B0(n3868), .B1(
        image_data[422]), .Y(n4024) );
  AOI22XL U5645 ( .A0(n3942), .A1(image_data[358]), .B0(n3943), .B1(
        image_data[486]), .Y(n4023) );
  AOI22XL U5646 ( .A0(n3865), .A1(image_data[326]), .B0(n3941), .B1(
        image_data[454]), .Y(n4025) );
  AOI22XL U5647 ( .A0(n3867), .A1(image_data[262]), .B0(n3866), .B1(
        image_data[390]), .Y(n4026) );
  NAND4XL U5648 ( .A(n4058), .B(n4057), .C(n4056), .D(n4055), .Y(n4059) );
  AOI22XL U5649 ( .A0(n3897), .A1(image_data[62]), .B0(n3896), .B1(
        image_data[190]), .Y(n4056) );
  AOI22XL U5650 ( .A0(n3928), .A1(image_data[94]), .B0(n3929), .B1(
        image_data[222]), .Y(n4057) );
  AOI22XL U5651 ( .A0(n3894), .A1(image_data[30]), .B0(n3893), .B1(
        image_data[158]), .Y(n4058) );
  NAND4XL U5652 ( .A(n4054), .B(n4053), .C(n4052), .D(n4051), .Y(n4060) );
  AOI22XL U5653 ( .A0(n3886), .A1(image_data[14]), .B0(n3885), .B1(
        image_data[142]), .Y(n4054) );
  AOI22XL U5654 ( .A0(n3887), .A1(image_data[110]), .B0(n3936), .B1(
        image_data[238]), .Y(n4051) );
  AOI22XL U5655 ( .A0(n4708), .A1(image_data[78]), .B0(n3934), .B1(
        image_data[206]), .Y(n4053) );
  NAND4XL U5656 ( .A(n4050), .B(n4049), .C(n4048), .D(n4047), .Y(n4061) );
  AOI22XL U5657 ( .A0(n3876), .A1(image_data[22]), .B0(n3875), .B1(
        image_data[150]), .Y(n4050) );
  AOI22XL U5658 ( .A0(n4722), .A1(image_data[118]), .B0(n3949), .B1(
        image_data[246]), .Y(n4047) );
  AOI22XL U5659 ( .A0(n4720), .A1(image_data[86]), .B0(n3948), .B1(
        image_data[214]), .Y(n4049) );
  NAND4XL U5660 ( .A(n4046), .B(n4045), .C(n4044), .D(n4043), .Y(n4062) );
  AOI22XL U5661 ( .A0(n3867), .A1(image_data[6]), .B0(n3866), .B1(
        image_data[134]), .Y(n4046) );
  AOI22XL U5662 ( .A0(n3865), .A1(image_data[70]), .B0(n3941), .B1(
        image_data[198]), .Y(n4045) );
  AOI22XL U5663 ( .A0(n3942), .A1(image_data[102]), .B0(n3943), .B1(
        image_data[230]), .Y(n4043) );
  NAND4XL U5664 ( .A(n4038), .B(n4037), .C(n4036), .D(n4035), .Y(n4039) );
  AOI22XL U5665 ( .A0(n3897), .A1(image_data[318]), .B0(n3896), .B1(
        image_data[446]), .Y(n4036) );
  AOI22XL U5666 ( .A0(n3791), .A1(image_data[350]), .B0(n3929), .B1(
        image_data[478]), .Y(n4037) );
  AOI22XL U5667 ( .A0(n3894), .A1(image_data[286]), .B0(n3893), .B1(
        image_data[414]), .Y(n4038) );
  NAND4XL U5668 ( .A(n4034), .B(n4033), .C(n4032), .D(n4031), .Y(n4040) );
  AOI22XL U5669 ( .A0(n3886), .A1(image_data[270]), .B0(n3885), .B1(
        image_data[398]), .Y(n4034) );
  AOI22XL U5670 ( .A0(n3887), .A1(image_data[366]), .B0(n3936), .B1(
        image_data[494]), .Y(n4031) );
  AOI22XL U5671 ( .A0(n4708), .A1(image_data[334]), .B0(n3934), .B1(
        image_data[462]), .Y(n4033) );
  NAND4XL U5672 ( .A(n4030), .B(n4029), .C(n4028), .D(n4027), .Y(n4041) );
  AOI22XL U5673 ( .A0(n3876), .A1(image_data[278]), .B0(n3875), .B1(
        image_data[406]), .Y(n4030) );
  AOI22XL U5674 ( .A0(n4722), .A1(image_data[374]), .B0(n3949), .B1(
        image_data[502]), .Y(n4027) );
  AOI22XL U5675 ( .A0(n4720), .A1(image_data[342]), .B0(n3948), .B1(
        image_data[470]), .Y(n4029) );
  NAND2XL U5676 ( .A(n5809), .B(op2[2]), .Y(n6800) );
  INVXL U5677 ( .A(n6123), .Y(n6029) );
  NAND4XL U5678 ( .A(n4088), .B(n4087), .C(n4086), .D(n4085), .Y(n4104) );
  AOI22XL U5679 ( .A0(n3897), .A1(image_data[67]), .B0(n3896), .B1(
        image_data[195]), .Y(n4087) );
  AOI22XL U5680 ( .A0(n3928), .A1(image_data[99]), .B0(n3929), .B1(
        image_data[227]), .Y(n4085) );
  AOI22XL U5681 ( .A0(n3894), .A1(image_data[35]), .B0(n3893), .B1(
        image_data[163]), .Y(n4086) );
  NAND4XL U5682 ( .A(n4100), .B(n4099), .C(n4098), .D(n4097), .Y(n4101) );
  AOI22XL U5683 ( .A0(n3876), .A1(image_data[27]), .B0(n3875), .B1(
        image_data[155]), .Y(n4100) );
  AOI22XL U5684 ( .A0(n3879), .A1(image_data[59]), .B0(n3878), .B1(
        image_data[187]), .Y(n4098) );
  AOI22XL U5685 ( .A0(n3877), .A1(image_data[123]), .B0(n3949), .B1(
        image_data[251]), .Y(n4097) );
  NAND4XL U5686 ( .A(n4096), .B(n4095), .C(n4094), .D(n4093), .Y(n4102) );
  AOI22XL U5687 ( .A0(n3867), .A1(image_data[11]), .B0(n3866), .B1(
        image_data[139]), .Y(n4096) );
  AOI22XL U5688 ( .A0(n4753), .A1(image_data[75]), .B0(n3941), .B1(
        image_data[203]), .Y(n4095) );
  AOI22XL U5689 ( .A0(n3942), .A1(image_data[107]), .B0(n3943), .B1(
        image_data[235]), .Y(n4093) );
  NAND4XL U5690 ( .A(n4092), .B(n4091), .C(n4090), .D(n4089), .Y(n4103) );
  AOI22XL U5691 ( .A0(n3888), .A1(image_data[51]), .B0(n4763), .B1(
        image_data[179]), .Y(n4090) );
  AOI22XL U5692 ( .A0(n3886), .A1(image_data[19]), .B0(n3885), .B1(
        image_data[147]), .Y(n4092) );
  AOI22XL U5693 ( .A0(n3887), .A1(image_data[115]), .B0(n3936), .B1(
        image_data[243]), .Y(n4089) );
  NAND4XL U5694 ( .A(n4068), .B(n4067), .C(n4066), .D(n4065), .Y(n4084) );
  AOI22XL U5695 ( .A0(n3894), .A1(image_data[291]), .B0(n4702), .B1(
        image_data[419]), .Y(n4066) );
  AOI22XL U5696 ( .A0(n3897), .A1(image_data[323]), .B0(n3896), .B1(
        image_data[451]), .Y(n4067) );
  AOI22XL U5697 ( .A0(n3928), .A1(image_data[355]), .B0(n3929), .B1(
        image_data[483]), .Y(n4065) );
  NAND4XL U5698 ( .A(n4080), .B(n4079), .C(n4078), .D(n4077), .Y(n4081) );
  AOI22XL U5699 ( .A0(n3876), .A1(image_data[283]), .B0(n3875), .B1(
        image_data[411]), .Y(n4080) );
  AOI22XL U5700 ( .A0(n3879), .A1(image_data[315]), .B0(n3878), .B1(
        image_data[443]), .Y(n4078) );
  AOI22XL U5701 ( .A0(n3877), .A1(image_data[379]), .B0(n3949), .B1(
        image_data[507]), .Y(n4077) );
  NAND4XL U5702 ( .A(n4076), .B(n4075), .C(n4074), .D(n4073), .Y(n4082) );
  AOI22XL U5703 ( .A0(n3867), .A1(image_data[267]), .B0(n3866), .B1(
        image_data[395]), .Y(n4076) );
  AOI22XL U5704 ( .A0(n3865), .A1(image_data[331]), .B0(n3941), .B1(
        image_data[459]), .Y(n4075) );
  AOI22XL U5705 ( .A0(n3869), .A1(image_data[299]), .B0(n3868), .B1(
        image_data[427]), .Y(n4074) );
  NAND4XL U5706 ( .A(n4072), .B(n4071), .C(n4070), .D(n4069), .Y(n4083) );
  AOI22XL U5707 ( .A0(n3886), .A1(image_data[275]), .B0(n4707), .B1(
        image_data[403]), .Y(n4072) );
  AOI22XL U5708 ( .A0(n3887), .A1(image_data[371]), .B0(n3936), .B1(
        image_data[499]), .Y(n4069) );
  AOI22XL U5709 ( .A0(n3888), .A1(image_data[307]), .B0(n3935), .B1(
        image_data[435]), .Y(n4070) );
  AOI22XL U5710 ( .A0(n3935), .A1(image_data[364]), .B0(n3888), .B1(
        image_data[492]), .Y(n4242) );
  AOI22XL U5711 ( .A0(n3887), .A1(image_data[300]), .B0(n3936), .B1(
        image_data[428]), .Y(n4243) );
  AOI22XL U5712 ( .A0(n3884), .A1(image_data[268]), .B0(n3934), .B1(
        image_data[396]), .Y(n4245) );
  AOI22XL U5713 ( .A0(n4707), .A1(image_data[332]), .B0(n3886), .B1(
        image_data[460]), .Y(n4244) );
  NAND4XL U5714 ( .A(n4269), .B(n4268), .C(n4267), .D(n4266), .Y(n4270) );
  AOI22XL U5715 ( .A0(n3928), .A1(image_data[28]), .B0(n3929), .B1(
        image_data[156]), .Y(n4269) );
  AOI22XL U5716 ( .A0(n3896), .A1(image_data[124]), .B0(n3897), .B1(
        image_data[252]), .Y(n4266) );
  AOI22XL U5717 ( .A0(n3893), .A1(image_data[92]), .B0(n3894), .B1(
        image_data[220]), .Y(n4268) );
  NAND4XL U5718 ( .A(n4261), .B(n4260), .C(n4259), .D(n4258), .Y(n4272) );
  AOI22XL U5719 ( .A0(n4719), .A1(image_data[84]), .B0(n3876), .B1(
        image_data[212]), .Y(n4260) );
  AOI22XL U5720 ( .A0(n3877), .A1(image_data[52]), .B0(n3949), .B1(
        image_data[180]), .Y(n4259) );
  AOI22XL U5721 ( .A0(n3874), .A1(image_data[20]), .B0(n3948), .B1(
        image_data[148]), .Y(n4261) );
  NAND4XL U5722 ( .A(n4257), .B(n4256), .C(n4255), .D(n4254), .Y(n4273) );
  AOI22XL U5723 ( .A0(n3866), .A1(image_data[68]), .B0(n3867), .B1(
        image_data[196]), .Y(n4256) );
  AOI22XL U5724 ( .A0(n3865), .A1(image_data[4]), .B0(n3941), .B1(
        image_data[132]), .Y(n4257) );
  AOI22XL U5725 ( .A0(n3942), .A1(image_data[36]), .B0(n3943), .B1(
        image_data[164]), .Y(n4255) );
  NAND4XL U5726 ( .A(n4265), .B(n4264), .C(n4263), .D(n4262), .Y(n4271) );
  AOI22XL U5727 ( .A0(n4707), .A1(image_data[76]), .B0(n3886), .B1(
        image_data[204]), .Y(n4264) );
  AOI22XL U5728 ( .A0(n3884), .A1(image_data[12]), .B0(n3934), .B1(
        image_data[140]), .Y(n4265) );
  AOI22XL U5729 ( .A0(n3887), .A1(image_data[44]), .B0(n3936), .B1(
        image_data[172]), .Y(n4263) );
  NAND4XL U5730 ( .A(n4249), .B(n4248), .C(n4247), .D(n4246), .Y(n4250) );
  AOI22XL U5731 ( .A0(n3896), .A1(image_data[380]), .B0(n3897), .B1(
        image_data[508]), .Y(n4246) );
  AOI22XL U5732 ( .A0(n3928), .A1(image_data[284]), .B0(n3929), .B1(
        image_data[412]), .Y(n4249) );
  AOI22XL U5733 ( .A0(n3893), .A1(image_data[348]), .B0(n3894), .B1(
        image_data[476]), .Y(n4248) );
  NAND4XL U5734 ( .A(n4241), .B(n4240), .C(n4239), .D(n4238), .Y(n4252) );
  AOI22XL U5735 ( .A0(n4719), .A1(image_data[340]), .B0(n3876), .B1(
        image_data[468]), .Y(n4240) );
  AOI22XL U5736 ( .A0(n3877), .A1(image_data[308]), .B0(n3949), .B1(
        image_data[436]), .Y(n4239) );
  AOI22XL U5737 ( .A0(n3874), .A1(image_data[276]), .B0(n3948), .B1(
        image_data[404]), .Y(n4241) );
  NAND4XL U5738 ( .A(n4237), .B(n4236), .C(n4235), .D(n4234), .Y(n4253) );
  AOI22XL U5739 ( .A0(n3866), .A1(image_data[324]), .B0(n3867), .B1(
        image_data[452]), .Y(n4236) );
  AOI22XL U5740 ( .A0(n3865), .A1(image_data[260]), .B0(n3941), .B1(
        image_data[388]), .Y(n4237) );
  AOI22XL U5741 ( .A0(n3942), .A1(image_data[292]), .B0(n3943), .B1(
        image_data[420]), .Y(n4235) );
  AOI22XL U5742 ( .A0(n3884), .A1(image_data[340]), .B0(n3934), .B1(
        image_data[468]), .Y(n4156) );
  AOI22XL U5743 ( .A0(n3887), .A1(image_data[372]), .B0(n3936), .B1(
        image_data[500]), .Y(n4154) );
  AOI22XL U5744 ( .A0(n3888), .A1(image_data[308]), .B0(n4763), .B1(
        image_data[436]), .Y(n4155) );
  AOI22XL U5745 ( .A0(n3886), .A1(image_data[276]), .B0(n3885), .B1(
        image_data[404]), .Y(n4157) );
  NAND4XL U5746 ( .A(n4185), .B(n4184), .C(n4183), .D(n4182), .Y(n4186) );
  AOI22XL U5747 ( .A0(n3876), .A1(image_data[28]), .B0(n3875), .B1(
        image_data[156]), .Y(n4185) );
  AOI22XL U5748 ( .A0(n3877), .A1(image_data[124]), .B0(n3949), .B1(
        image_data[252]), .Y(n4182) );
  AOI22XL U5749 ( .A0(n3874), .A1(image_data[92]), .B0(n3948), .B1(
        image_data[220]), .Y(n4184) );
  NAND4XL U5750 ( .A(n4181), .B(n4180), .C(n4179), .D(n4178), .Y(n4187) );
  AOI22XL U5751 ( .A0(n3867), .A1(image_data[12]), .B0(n3866), .B1(
        image_data[140]), .Y(n4181) );
  AOI22XL U5752 ( .A0(n3865), .A1(image_data[76]), .B0(n3941), .B1(
        image_data[204]), .Y(n4180) );
  AOI22XL U5753 ( .A0(n3942), .A1(image_data[108]), .B0(n3943), .B1(
        image_data[236]), .Y(n4178) );
  NAND4XL U5754 ( .A(n4173), .B(n4172), .C(n4171), .D(n4170), .Y(n4189) );
  AOI22XL U5755 ( .A0(n3364), .A1(image_data[4]), .B0(n4681), .B1(
        image_data[132]), .Y(n4173) );
  AOI22XL U5756 ( .A0(n3897), .A1(image_data[68]), .B0(n3896), .B1(
        image_data[196]), .Y(n4172) );
  AOI22XL U5757 ( .A0(n3928), .A1(image_data[100]), .B0(n3929), .B1(
        image_data[228]), .Y(n4170) );
  NAND4XL U5758 ( .A(n4177), .B(n4176), .C(n4175), .D(n4174), .Y(n4188) );
  AOI22XL U5759 ( .A0(n3886), .A1(image_data[20]), .B0(n3885), .B1(
        image_data[148]), .Y(n4177) );
  AOI22XL U5760 ( .A0(n3887), .A1(image_data[116]), .B0(n3936), .B1(
        image_data[244]), .Y(n4174) );
  AOI22XL U5761 ( .A0(n3884), .A1(image_data[84]), .B0(n3934), .B1(
        image_data[212]), .Y(n4176) );
  NAND4XL U5762 ( .A(n4165), .B(n4164), .C(n4163), .D(n4162), .Y(n4166) );
  AOI22XL U5763 ( .A0(n3876), .A1(image_data[284]), .B0(n3875), .B1(
        image_data[412]), .Y(n4165) );
  AOI22XL U5764 ( .A0(n3877), .A1(image_data[380]), .B0(n3949), .B1(
        image_data[508]), .Y(n4162) );
  AOI22XL U5765 ( .A0(n3874), .A1(image_data[348]), .B0(n3948), .B1(
        image_data[476]), .Y(n4164) );
  NAND4XL U5766 ( .A(n4161), .B(n4160), .C(n4159), .D(n4158), .Y(n4167) );
  AOI22XL U5767 ( .A0(n3867), .A1(image_data[268]), .B0(n3866), .B1(
        image_data[396]), .Y(n4161) );
  AOI22XL U5768 ( .A0(n3865), .A1(image_data[332]), .B0(n3941), .B1(
        image_data[460]), .Y(n4160) );
  AOI22XL U5769 ( .A0(n3942), .A1(image_data[364]), .B0(n3943), .B1(
        image_data[492]), .Y(n4158) );
  NAND4XL U5770 ( .A(n4153), .B(n4152), .C(n4151), .D(n4150), .Y(n4169) );
  AOI22XL U5771 ( .A0(n3364), .A1(image_data[260]), .B0(n4681), .B1(
        image_data[388]), .Y(n4153) );
  AOI22XL U5772 ( .A0(n3897), .A1(image_data[324]), .B0(n3896), .B1(
        image_data[452]), .Y(n4152) );
  AOI22XL U5773 ( .A0(n3928), .A1(image_data[356]), .B0(n3929), .B1(
        image_data[484]), .Y(n4150) );
  AOI22XL U5774 ( .A0(n3879), .A1(image_data[307]), .B0(n3878), .B1(
        image_data[435]), .Y(n4113) );
  AOI22XL U5775 ( .A0(n3874), .A1(image_data[339]), .B0(n3948), .B1(
        image_data[467]), .Y(n4114) );
  AOI22XL U5776 ( .A0(n3877), .A1(image_data[371]), .B0(n3949), .B1(
        image_data[499]), .Y(n4112) );
  AOI22XL U5777 ( .A0(n3876), .A1(image_data[275]), .B0(n3875), .B1(
        image_data[403]), .Y(n4115) );
  NAND4XL U5778 ( .A(n4143), .B(n4142), .C(n4141), .D(n4140), .Y(n4144) );
  AOI22XL U5779 ( .A0(n3897), .A1(image_data[59]), .B0(n3896), .B1(
        image_data[187]), .Y(n4141) );
  AOI22XL U5780 ( .A0(n3928), .A1(image_data[91]), .B0(n3929), .B1(
        image_data[219]), .Y(n4142) );
  AOI22XL U5781 ( .A0(n3894), .A1(image_data[27]), .B0(n3893), .B1(
        image_data[155]), .Y(n4143) );
  NAND4XL U5782 ( .A(n4139), .B(n4138), .C(n4137), .D(n4136), .Y(n4145) );
  AOI22XL U5783 ( .A0(n3886), .A1(image_data[11]), .B0(n3885), .B1(
        image_data[139]), .Y(n4139) );
  AOI22XL U5784 ( .A0(n3887), .A1(image_data[107]), .B0(n3936), .B1(
        image_data[235]), .Y(n4136) );
  AOI22XL U5785 ( .A0(n3884), .A1(image_data[75]), .B0(n3934), .B1(
        image_data[203]), .Y(n4138) );
  NAND4XL U5786 ( .A(n4131), .B(n4130), .C(n4129), .D(n4128), .Y(n4147) );
  AOI22XL U5787 ( .A0(n3867), .A1(image_data[3]), .B0(n3866), .B1(
        image_data[131]), .Y(n4131) );
  AOI22XL U5788 ( .A0(n3865), .A1(image_data[67]), .B0(n3941), .B1(
        image_data[195]), .Y(n4130) );
  AOI22XL U5789 ( .A0(n3942), .A1(image_data[99]), .B0(n3943), .B1(
        image_data[227]), .Y(n4128) );
  NAND4XL U5790 ( .A(n4135), .B(n4134), .C(n4133), .D(n4132), .Y(n4146) );
  AOI22XL U5791 ( .A0(n3876), .A1(image_data[19]), .B0(n3875), .B1(
        image_data[147]), .Y(n4135) );
  AOI22XL U5792 ( .A0(n3877), .A1(image_data[115]), .B0(n3949), .B1(
        image_data[243]), .Y(n4132) );
  AOI22XL U5793 ( .A0(n3874), .A1(image_data[83]), .B0(n3948), .B1(
        image_data[211]), .Y(n4134) );
  NAND4XL U5794 ( .A(n4123), .B(n4122), .C(n4121), .D(n4120), .Y(n4124) );
  AOI22XL U5795 ( .A0(n3897), .A1(image_data[315]), .B0(n3896), .B1(
        image_data[443]), .Y(n4121) );
  AOI22XL U5796 ( .A0(n3928), .A1(image_data[347]), .B0(n3929), .B1(
        image_data[475]), .Y(n4122) );
  AOI22XL U5797 ( .A0(n3894), .A1(image_data[283]), .B0(n3893), .B1(
        image_data[411]), .Y(n4123) );
  NAND4XL U5798 ( .A(n4119), .B(n4118), .C(n4117), .D(n4116), .Y(n4125) );
  AOI22XL U5799 ( .A0(n3886), .A1(image_data[267]), .B0(n3885), .B1(
        image_data[395]), .Y(n4119) );
  AOI22XL U5800 ( .A0(n3887), .A1(image_data[363]), .B0(n3936), .B1(
        image_data[491]), .Y(n4116) );
  AOI22XL U5801 ( .A0(n3884), .A1(image_data[331]), .B0(n3934), .B1(
        image_data[459]), .Y(n4118) );
  NAND4XL U5802 ( .A(n4111), .B(n4110), .C(n4109), .D(n4108), .Y(n4127) );
  AOI22XL U5803 ( .A0(n3867), .A1(image_data[259]), .B0(n3866), .B1(
        image_data[387]), .Y(n4111) );
  AOI22XL U5804 ( .A0(n4753), .A1(image_data[323]), .B0(n3941), .B1(
        image_data[451]), .Y(n4110) );
  AOI22XL U5805 ( .A0(n4754), .A1(image_data[355]), .B0(n3943), .B1(
        image_data[483]), .Y(n4108) );
  AOI22XL U5806 ( .A0(n3886), .A1(image_data[277]), .B0(n3885), .B1(
        image_data[405]), .Y(n3988) );
  NAND4XL U5807 ( .A(n3721), .B(n3720), .C(n3719), .D(n3718), .Y(n3722) );
  AOI22XL U5808 ( .A0(n3876), .A1(image_data[30]), .B0(n3875), .B1(
        image_data[158]), .Y(n3721) );
  AOI22XL U5809 ( .A0(n3879), .A1(image_data[62]), .B0(n3878), .B1(
        image_data[190]), .Y(n3719) );
  AOI22XL U5810 ( .A0(n3877), .A1(image_data[126]), .B0(n3949), .B1(
        image_data[254]), .Y(n3718) );
  NAND4XL U5811 ( .A(n3717), .B(n3716), .C(n3715), .D(n3714), .Y(n3723) );
  AOI22XL U5812 ( .A0(n3867), .A1(image_data[14]), .B0(n3866), .B1(
        image_data[142]), .Y(n3717) );
  AOI22XL U5813 ( .A0(n4753), .A1(image_data[78]), .B0(n3941), .B1(
        image_data[206]), .Y(n3716) );
  AOI22XL U5814 ( .A0(n3869), .A1(image_data[46]), .B0(n3868), .B1(
        image_data[174]), .Y(n3715) );
  NAND4XL U5815 ( .A(n3709), .B(n3708), .C(n3707), .D(n3706), .Y(n3725) );
  AOI22XL U5816 ( .A0(n3364), .A1(image_data[6]), .B0(n4681), .B1(
        image_data[134]), .Y(n3709) );
  AOI22XL U5817 ( .A0(n3897), .A1(image_data[70]), .B0(n3896), .B1(
        image_data[198]), .Y(n3708) );
  AOI22XL U5818 ( .A0(n3928), .A1(image_data[102]), .B0(n3929), .B1(
        image_data[230]), .Y(n3706) );
  NAND4XL U5819 ( .A(n3713), .B(n3712), .C(n3711), .D(n3710), .Y(n3724) );
  AOI22XL U5820 ( .A0(n3888), .A1(image_data[54]), .B0(n4763), .B1(
        image_data[182]), .Y(n3711) );
  AOI22XL U5821 ( .A0(n3886), .A1(image_data[22]), .B0(n3885), .B1(
        image_data[150]), .Y(n3713) );
  AOI22XL U5822 ( .A0(n3887), .A1(image_data[118]), .B0(n3936), .B1(
        image_data[246]), .Y(n3710) );
  NAND4XL U5823 ( .A(n3701), .B(n3700), .C(n3699), .D(n3698), .Y(n3702) );
  AOI22XL U5824 ( .A0(n3876), .A1(image_data[286]), .B0(n3875), .B1(
        image_data[414]), .Y(n3701) );
  AOI22XL U5825 ( .A0(n3879), .A1(image_data[318]), .B0(n3878), .B1(
        image_data[446]), .Y(n3699) );
  AOI22XL U5826 ( .A0(n3877), .A1(image_data[382]), .B0(n3949), .B1(
        image_data[510]), .Y(n3698) );
  NAND4XL U5827 ( .A(n3697), .B(n3696), .C(n3695), .D(n3694), .Y(n3703) );
  AOI22XL U5828 ( .A0(n3867), .A1(image_data[270]), .B0(n3866), .B1(
        image_data[398]), .Y(n3697) );
  AOI22XL U5829 ( .A0(n4753), .A1(image_data[334]), .B0(n3941), .B1(
        image_data[462]), .Y(n3696) );
  AOI22XL U5830 ( .A0(n3869), .A1(image_data[302]), .B0(n3868), .B1(
        image_data[430]), .Y(n3695) );
  NAND4XL U5831 ( .A(n3689), .B(n3688), .C(n3687), .D(n3686), .Y(n3705) );
  AOI22XL U5832 ( .A0(n3364), .A1(image_data[262]), .B0(n4681), .B1(
        image_data[390]), .Y(n3689) );
  AOI22XL U5833 ( .A0(n3897), .A1(image_data[326]), .B0(n3896), .B1(
        image_data[454]), .Y(n3688) );
  AOI22XL U5834 ( .A0(n3928), .A1(image_data[358]), .B0(n3929), .B1(
        image_data[486]), .Y(n3686) );
  NAND4XL U5835 ( .A(n3693), .B(n3692), .C(n3691), .D(n3690), .Y(n3704) );
  AOI22XL U5836 ( .A0(n3888), .A1(image_data[310]), .B0(n4763), .B1(
        image_data[438]), .Y(n3691) );
  AOI22XL U5837 ( .A0(n3886), .A1(image_data[278]), .B0(n3885), .B1(
        image_data[406]), .Y(n3693) );
  AOI22XL U5838 ( .A0(n3887), .A1(image_data[374]), .B0(n3936), .B1(
        image_data[502]), .Y(n3690) );
  AOI22XL U5839 ( .A0(n3935), .A1(image_data[375]), .B0(n3888), .B1(
        image_data[503]), .Y(n3564) );
  AOI22XL U5840 ( .A0(n3887), .A1(image_data[311]), .B0(n3936), .B1(
        image_data[439]), .Y(n3565) );
  AOI22XL U5841 ( .A0(n3884), .A1(image_data[279]), .B0(n3934), .B1(
        image_data[407]), .Y(n3567) );
  AOI22XL U5842 ( .A0(n3885), .A1(image_data[343]), .B0(n3886), .B1(
        image_data[471]), .Y(n3566) );
  NAND4XL U5843 ( .A(n3595), .B(n3594), .C(n3593), .D(n3592), .Y(n3596) );
  AOI22XL U5844 ( .A0(n3875), .A1(image_data[95]), .B0(n3876), .B1(
        image_data[223]), .Y(n3594) );
  AOI22XL U5845 ( .A0(n3877), .A1(image_data[63]), .B0(n3949), .B1(
        image_data[191]), .Y(n3593) );
  AOI22XL U5846 ( .A0(n3874), .A1(image_data[31]), .B0(n3948), .B1(
        image_data[159]), .Y(n3595) );
  NAND4XL U5847 ( .A(n3591), .B(n3590), .C(n3589), .D(n3588), .Y(n3597) );
  AOI22XL U5848 ( .A0(n3866), .A1(image_data[79]), .B0(n3867), .B1(
        image_data[207]), .Y(n3590) );
  AOI22XL U5849 ( .A0(n3865), .A1(image_data[15]), .B0(n3941), .B1(
        image_data[143]), .Y(n3591) );
  AOI22XL U5850 ( .A0(n3942), .A1(image_data[47]), .B0(n3943), .B1(
        image_data[175]), .Y(n3589) );
  NAND4XL U5851 ( .A(n3583), .B(n3582), .C(n3581), .D(n3580), .Y(n3599) );
  AOI22XL U5852 ( .A0(n4681), .A1(image_data[71]), .B0(n3364), .B1(
        image_data[199]), .Y(n3582) );
  AOI22XL U5853 ( .A0(n3897), .A1(image_data[7]), .B0(n3896), .B1(
        image_data[135]), .Y(n3583) );
  AOI22XL U5854 ( .A0(n3928), .A1(image_data[39]), .B0(n3929), .B1(
        image_data[167]), .Y(n3581) );
  NAND4XL U5855 ( .A(n3587), .B(n3586), .C(n3585), .D(n3584), .Y(n3598) );
  AOI22XL U5856 ( .A0(n3885), .A1(image_data[87]), .B0(n3886), .B1(
        image_data[215]), .Y(n3586) );
  AOI22XL U5857 ( .A0(n3884), .A1(image_data[23]), .B0(n3934), .B1(
        image_data[151]), .Y(n3587) );
  AOI22XL U5858 ( .A0(n3887), .A1(image_data[55]), .B0(n3936), .B1(
        image_data[183]), .Y(n3585) );
  NAND4XL U5859 ( .A(n3575), .B(n3574), .C(n3573), .D(n3572), .Y(n3576) );
  AOI22XL U5860 ( .A0(n3875), .A1(image_data[351]), .B0(n3876), .B1(
        image_data[479]), .Y(n3574) );
  AOI22XL U5861 ( .A0(n3877), .A1(image_data[319]), .B0(n3949), .B1(
        image_data[447]), .Y(n3573) );
  AOI22XL U5862 ( .A0(n3874), .A1(image_data[287]), .B0(n3948), .B1(
        image_data[415]), .Y(n3575) );
  NAND4XL U5863 ( .A(n3571), .B(n3570), .C(n3569), .D(n3568), .Y(n3577) );
  AOI22XL U5864 ( .A0(n3865), .A1(image_data[271]), .B0(n4433), .B1(
        image_data[399]), .Y(n3571) );
  AOI22XL U5865 ( .A0(n3866), .A1(image_data[335]), .B0(n3867), .B1(
        image_data[463]), .Y(n3570) );
  AOI22XL U5866 ( .A0(n3942), .A1(image_data[303]), .B0(n3943), .B1(
        image_data[431]), .Y(n3569) );
  NAND4XL U5867 ( .A(n3563), .B(n3562), .C(n3561), .D(n3560), .Y(n3579) );
  AOI22XL U5868 ( .A0(n3791), .A1(image_data[295]), .B0(n3929), .B1(
        image_data[423]), .Y(n3561) );
  AOI22XL U5869 ( .A0(n3897), .A1(image_data[263]), .B0(n3896), .B1(
        image_data[391]), .Y(n3563) );
  AOI22XL U5870 ( .A0(n3895), .A1(image_data[327]), .B0(n3364), .B1(
        image_data[455]), .Y(n3562) );
  AOI22XL U5871 ( .A0(n3869), .A1(image_data[295]), .B0(n3868), .B1(
        image_data[423]), .Y(n3603) );
  AOI22XL U5872 ( .A0(n3942), .A1(image_data[359]), .B0(n3943), .B1(
        image_data[487]), .Y(n3602) );
  AOI22XL U5873 ( .A0(n3865), .A1(image_data[327]), .B0(n3941), .B1(
        image_data[455]), .Y(n3604) );
  AOI22XL U5874 ( .A0(n3867), .A1(image_data[263]), .B0(n3866), .B1(
        image_data[391]), .Y(n3605) );
  NAND4XL U5875 ( .A(n3637), .B(n3636), .C(n3635), .D(n3634), .Y(n3638) );
  AOI22XL U5876 ( .A0(n3897), .A1(image_data[63]), .B0(n3896), .B1(
        image_data[191]), .Y(n3635) );
  AOI22XL U5877 ( .A0(n3791), .A1(image_data[95]), .B0(n3929), .B1(
        image_data[223]), .Y(n3636) );
  AOI22XL U5878 ( .A0(n3894), .A1(image_data[31]), .B0(n3893), .B1(
        image_data[159]), .Y(n3637) );
  NAND4XL U5879 ( .A(n3633), .B(n3632), .C(n3631), .D(n3630), .Y(n3639) );
  AOI22XL U5880 ( .A0(n3886), .A1(image_data[15]), .B0(n3885), .B1(
        image_data[143]), .Y(n3633) );
  AOI22XL U5881 ( .A0(n3887), .A1(image_data[111]), .B0(n3936), .B1(
        image_data[239]), .Y(n3630) );
  AOI22XL U5882 ( .A0(n4708), .A1(image_data[79]), .B0(n3934), .B1(
        image_data[207]), .Y(n3632) );
  NAND4XL U5883 ( .A(n3629), .B(n3628), .C(n3627), .D(n3626), .Y(n3640) );
  AOI22XL U5884 ( .A0(n3876), .A1(image_data[23]), .B0(n3875), .B1(
        image_data[151]), .Y(n3629) );
  AOI22XL U5885 ( .A0(n4722), .A1(image_data[119]), .B0(n3949), .B1(
        image_data[247]), .Y(n3626) );
  AOI22XL U5886 ( .A0(n4720), .A1(image_data[87]), .B0(n3948), .B1(
        image_data[215]), .Y(n3628) );
  NAND4XL U5887 ( .A(n3625), .B(n3624), .C(n3623), .D(n3622), .Y(n3641) );
  AOI22XL U5888 ( .A0(n3867), .A1(image_data[7]), .B0(n3866), .B1(
        image_data[135]), .Y(n3625) );
  AOI22XL U5889 ( .A0(n3865), .A1(image_data[71]), .B0(n3941), .B1(
        image_data[199]), .Y(n3624) );
  AOI22XL U5890 ( .A0(n3942), .A1(image_data[103]), .B0(n3943), .B1(
        image_data[231]), .Y(n3622) );
  NAND4XL U5891 ( .A(n3617), .B(n3616), .C(n3615), .D(n3614), .Y(n3618) );
  AOI22XL U5892 ( .A0(n4681), .A1(image_data[383]), .B0(n3364), .B1(
        image_data[511]), .Y(n3614) );
  AOI22XL U5893 ( .A0(n3897), .A1(image_data[319]), .B0(n3896), .B1(
        image_data[447]), .Y(n3615) );
  AOI22XL U5894 ( .A0(n3791), .A1(image_data[351]), .B0(n3929), .B1(
        image_data[479]), .Y(n3616) );
  NAND4XL U5895 ( .A(n3613), .B(n3612), .C(n3611), .D(n3610), .Y(n3619) );
  AOI22XL U5896 ( .A0(n3886), .A1(image_data[271]), .B0(n3885), .B1(
        image_data[399]), .Y(n3613) );
  AOI22XL U5897 ( .A0(n3887), .A1(image_data[367]), .B0(n3936), .B1(
        image_data[495]), .Y(n3610) );
  AOI22XL U5898 ( .A0(n4708), .A1(image_data[335]), .B0(n3934), .B1(
        image_data[463]), .Y(n3612) );
  NAND4XL U5899 ( .A(n3609), .B(n3608), .C(n3607), .D(n3606), .Y(n3620) );
  AOI22XL U5900 ( .A0(n3876), .A1(image_data[279]), .B0(n3875), .B1(
        image_data[407]), .Y(n3609) );
  AOI22XL U5901 ( .A0(n4722), .A1(image_data[375]), .B0(n3949), .B1(
        image_data[503]), .Y(n3606) );
  AOI22XL U5902 ( .A0(n4720), .A1(image_data[343]), .B0(n3948), .B1(
        image_data[471]), .Y(n3608) );
  NOR3XL U5903 ( .A(n8530), .B(n8528), .C(n6902), .Y(n6819) );
  NAND4XL U5904 ( .A(n3961), .B(n3960), .C(n3959), .D(n3958), .Y(n3977) );
  AOI22XL U5905 ( .A0(n3894), .A1(image_data[34]), .B0(n4702), .B1(
        image_data[162]), .Y(n3959) );
  AOI22XL U5906 ( .A0(n3897), .A1(image_data[66]), .B0(n3896), .B1(
        image_data[194]), .Y(n3960) );
  AOI22XL U5907 ( .A0(n3928), .A1(image_data[98]), .B0(n3929), .B1(
        image_data[226]), .Y(n3958) );
  NAND4XL U5908 ( .A(n3973), .B(n3972), .C(n3971), .D(n3970), .Y(n3974) );
  AOI22XL U5909 ( .A0(n3876), .A1(image_data[26]), .B0(n4719), .B1(
        image_data[154]), .Y(n3973) );
  AOI22XL U5910 ( .A0(n3879), .A1(image_data[58]), .B0(n4721), .B1(
        image_data[186]), .Y(n3971) );
  AOI22XL U5911 ( .A0(n3877), .A1(image_data[122]), .B0(n3949), .B1(
        image_data[250]), .Y(n3970) );
  NAND4XL U5912 ( .A(n3969), .B(n3968), .C(n3967), .D(n3966), .Y(n3975) );
  AOI22XL U5913 ( .A0(n3869), .A1(image_data[42]), .B0(n4714), .B1(
        image_data[170]), .Y(n3967) );
  AOI22XL U5914 ( .A0(n3867), .A1(image_data[10]), .B0(n3866), .B1(
        image_data[138]), .Y(n3969) );
  AOI22XL U5915 ( .A0(n3865), .A1(image_data[74]), .B0(n3941), .B1(
        image_data[202]), .Y(n3968) );
  NAND4XL U5916 ( .A(n3965), .B(n3964), .C(n3963), .D(n3962), .Y(n3976) );
  AOI22XL U5917 ( .A0(n3886), .A1(image_data[18]), .B0(n4707), .B1(
        image_data[146]), .Y(n3965) );
  AOI22XL U5918 ( .A0(n3887), .A1(image_data[114]), .B0(n3936), .B1(
        image_data[242]), .Y(n3962) );
  AOI22XL U5919 ( .A0(n3888), .A1(image_data[50]), .B0(n3935), .B1(
        image_data[178]), .Y(n3963) );
  NAND4XL U5920 ( .A(n3953), .B(n3952), .C(n3951), .D(n3950), .Y(n3954) );
  AOI22XL U5921 ( .A0(n3876), .A1(image_data[282]), .B0(n4719), .B1(
        image_data[410]), .Y(n3953) );
  AOI22XL U5922 ( .A0(n3879), .A1(image_data[314]), .B0(n4721), .B1(
        image_data[442]), .Y(n3951) );
  AOI22XL U5923 ( .A0(n3877), .A1(image_data[378]), .B0(n3949), .B1(
        image_data[506]), .Y(n3950) );
  NAND4XL U5924 ( .A(n3947), .B(n3946), .C(n3945), .D(n3944), .Y(n3955) );
  AOI22XL U5925 ( .A0(n3869), .A1(image_data[298]), .B0(n4714), .B1(
        image_data[426]), .Y(n3945) );
  AOI22XL U5926 ( .A0(n3867), .A1(image_data[266]), .B0(n3866), .B1(
        image_data[394]), .Y(n3947) );
  AOI22XL U5927 ( .A0(n3865), .A1(image_data[330]), .B0(n3941), .B1(
        image_data[458]), .Y(n3946) );
  NAND4XL U5928 ( .A(n3940), .B(n3939), .C(n3938), .D(n3937), .Y(n3956) );
  AOI22XL U5929 ( .A0(n3886), .A1(image_data[274]), .B0(n4707), .B1(
        image_data[402]), .Y(n3940) );
  AOI22XL U5930 ( .A0(n3887), .A1(image_data[370]), .B0(n3936), .B1(
        image_data[498]), .Y(n3937) );
  AOI22XL U5931 ( .A0(n3888), .A1(image_data[306]), .B0(n3935), .B1(
        image_data[434]), .Y(n3938) );
  NAND4XL U5932 ( .A(n3933), .B(n3932), .C(n3931), .D(n3930), .Y(n3957) );
  AOI22XL U5933 ( .A0(n3894), .A1(image_data[290]), .B0(n4702), .B1(
        image_data[418]), .Y(n3931) );
  AOI22XL U5934 ( .A0(n3364), .A1(image_data[258]), .B0(n4681), .B1(
        image_data[386]), .Y(n3933) );
  AOI22XL U5935 ( .A0(n3897), .A1(image_data[322]), .B0(n3896), .B1(
        image_data[450]), .Y(n3932) );
  NOR4XL U5936 ( .A(n3748), .B(n3747), .C(n3746), .D(n3745), .Y(n3770) );
  NOR4XL U5937 ( .A(n3768), .B(n3767), .C(n3766), .D(n3765), .Y(n3769) );
  NAND4XL U5938 ( .A(n3736), .B(n3735), .C(n3734), .D(n3733), .Y(n3747) );
  INVX1 U5939 ( .A(n6136), .Y(n5013) );
  AOI22XL U5940 ( .A0(op4[5]), .A1(n3517), .B0(n3516), .B1(n8525), .Y(N2763)
         );
  AOI22XL U5941 ( .A0(n3866), .A1(image_data[327]), .B0(n3867), .B1(
        image_data[455]), .Y(n4362) );
  AOI22XL U5942 ( .A0(n3865), .A1(image_data[263]), .B0(n3941), .B1(
        image_data[391]), .Y(n4363) );
  AOI22XL U5943 ( .A0(n5582), .A1(image_data[24]), .B0(n5581), .B1(
        image_data[152]), .Y(n5518) );
  AOI22XL U5944 ( .A0(n5570), .A1(image_data[8]), .B0(n5569), .B1(
        image_data[136]), .Y(n5514) );
  AOI22XL U5945 ( .A0(n5558), .A1(image_data[16]), .B0(n5557), .B1(
        image_data[144]), .Y(n5510) );
  AOI22XL U5946 ( .A0(n5546), .A1(image_data[0]), .B0(n5545), .B1(
        image_data[128]), .Y(n5506) );
  AOI22XL U5947 ( .A0(n5582), .A1(image_data[280]), .B0(n5581), .B1(
        image_data[408]), .Y(n5498) );
  AOI22XL U5948 ( .A0(n5570), .A1(image_data[264]), .B0(n5569), .B1(
        image_data[392]), .Y(n5494) );
  AOI22XL U5949 ( .A0(n5558), .A1(image_data[272]), .B0(n5557), .B1(
        image_data[400]), .Y(n5490) );
  AOI22XL U5950 ( .A0(n5582), .A1(image_data[25]), .B0(n5581), .B1(
        image_data[153]), .Y(n5434) );
  AOI22XL U5951 ( .A0(n5570), .A1(image_data[9]), .B0(n5569), .B1(
        image_data[137]), .Y(n5430) );
  AOI22XL U5952 ( .A0(n5558), .A1(image_data[17]), .B0(n5557), .B1(
        image_data[145]), .Y(n5426) );
  AOI22XL U5953 ( .A0(n5546), .A1(image_data[1]), .B0(n5545), .B1(
        image_data[129]), .Y(n5422) );
  AOI22XL U5954 ( .A0(n5582), .A1(image_data[281]), .B0(n5581), .B1(
        image_data[409]), .Y(n5414) );
  AOI22XL U5955 ( .A0(n5570), .A1(image_data[265]), .B0(n5569), .B1(
        image_data[393]), .Y(n5410) );
  AOI22XL U5956 ( .A0(n5558), .A1(image_data[273]), .B0(n5557), .B1(
        image_data[401]), .Y(n5406) );
  AOI22XL U5957 ( .A0(n5582), .A1(image_data[26]), .B0(n5581), .B1(
        image_data[154]), .Y(n4580) );
  AOI22XL U5958 ( .A0(n5570), .A1(image_data[10]), .B0(n5569), .B1(
        image_data[138]), .Y(n4576) );
  AOI22XL U5959 ( .A0(n5558), .A1(image_data[18]), .B0(n5557), .B1(
        image_data[146]), .Y(n4572) );
  AOI22XL U5960 ( .A0(n5546), .A1(image_data[2]), .B0(n5545), .B1(
        image_data[130]), .Y(n4568) );
  AOI22XL U5961 ( .A0(n5582), .A1(image_data[282]), .B0(n5581), .B1(
        image_data[410]), .Y(n4560) );
  AOI22XL U5962 ( .A0(n5570), .A1(image_data[266]), .B0(n5569), .B1(
        image_data[394]), .Y(n4548) );
  AOI22XL U5963 ( .A0(n5558), .A1(image_data[274]), .B0(n5557), .B1(
        image_data[402]), .Y(n4544) );
  AOI22XL U5964 ( .A0(n5582), .A1(image_data[27]), .B0(n5581), .B1(
        image_data[155]), .Y(n5592) );
  AOI22XL U5965 ( .A0(n5570), .A1(image_data[11]), .B0(n5569), .B1(
        image_data[139]), .Y(n5580) );
  AOI22XL U5966 ( .A0(n5558), .A1(image_data[19]), .B0(n5557), .B1(
        image_data[147]), .Y(n5568) );
  AOI22XL U5967 ( .A0(n5546), .A1(image_data[3]), .B0(n5545), .B1(
        image_data[131]), .Y(n5556) );
  AOI22XL U5968 ( .A0(n5582), .A1(image_data[283]), .B0(n5581), .B1(
        image_data[411]), .Y(n5540) );
  AOI22XL U5969 ( .A0(n5570), .A1(image_data[267]), .B0(n5569), .B1(
        image_data[395]), .Y(n5536) );
  AOI22XL U5970 ( .A0(n5558), .A1(image_data[275]), .B0(n5557), .B1(
        image_data[403]), .Y(n5532) );
  AOI22XL U5971 ( .A0(n5582), .A1(image_data[28]), .B0(n5581), .B1(
        image_data[156]), .Y(n5476) );
  AOI22XL U5972 ( .A0(n5570), .A1(image_data[12]), .B0(n5569), .B1(
        image_data[140]), .Y(n5472) );
  AOI22XL U5973 ( .A0(n5558), .A1(image_data[20]), .B0(n5557), .B1(
        image_data[148]), .Y(n5468) );
  AOI22XL U5974 ( .A0(n5546), .A1(image_data[4]), .B0(n5545), .B1(
        image_data[132]), .Y(n5464) );
  AOI22XL U5975 ( .A0(n5582), .A1(image_data[284]), .B0(n5581), .B1(
        image_data[412]), .Y(n5456) );
  AOI22XL U5976 ( .A0(n5570), .A1(image_data[268]), .B0(n5569), .B1(
        image_data[396]), .Y(n5452) );
  AOI22XL U5977 ( .A0(n5558), .A1(image_data[276]), .B0(n5557), .B1(
        image_data[404]), .Y(n5448) );
  AOI22XL U5978 ( .A0(n5582), .A1(image_data[29]), .B0(n5581), .B1(
        image_data[157]), .Y(n5392) );
  AOI22XL U5979 ( .A0(n5570), .A1(image_data[13]), .B0(n5569), .B1(
        image_data[141]), .Y(n5388) );
  AOI22XL U5980 ( .A0(n5558), .A1(image_data[21]), .B0(n5557), .B1(
        image_data[149]), .Y(n5384) );
  AOI22XL U5981 ( .A0(n5546), .A1(image_data[5]), .B0(n5545), .B1(
        image_data[133]), .Y(n5380) );
  AOI22XL U5982 ( .A0(n5582), .A1(image_data[285]), .B0(n5581), .B1(
        image_data[413]), .Y(n5372) );
  AOI22XL U5983 ( .A0(n5570), .A1(image_data[269]), .B0(n5569), .B1(
        image_data[397]), .Y(n5368) );
  AOI22XL U5984 ( .A0(n5558), .A1(image_data[277]), .B0(n5557), .B1(
        image_data[405]), .Y(n5364) );
  AOI22XL U5985 ( .A0(n5582), .A1(image_data[30]), .B0(n5581), .B1(
        image_data[158]), .Y(n5350) );
  AOI22XL U5986 ( .A0(n5570), .A1(image_data[14]), .B0(n5569), .B1(
        image_data[142]), .Y(n5346) );
  AOI22XL U5987 ( .A0(n5558), .A1(image_data[22]), .B0(n5557), .B1(
        image_data[150]), .Y(n5342) );
  AOI22XL U5988 ( .A0(n5546), .A1(image_data[6]), .B0(n5545), .B1(
        image_data[134]), .Y(n5338) );
  AOI22XL U5989 ( .A0(n5582), .A1(image_data[286]), .B0(n5581), .B1(
        image_data[414]), .Y(n5330) );
  AOI22XL U5990 ( .A0(n5570), .A1(image_data[270]), .B0(n5569), .B1(
        image_data[398]), .Y(n5326) );
  AOI22XL U5991 ( .A0(n5558), .A1(image_data[278]), .B0(n5557), .B1(
        image_data[406]), .Y(n5322) );
  AOI22XL U5992 ( .A0(n5582), .A1(image_data[31]), .B0(n5581), .B1(
        image_data[159]), .Y(n5308) );
  AOI22XL U5993 ( .A0(n5570), .A1(image_data[15]), .B0(n5569), .B1(
        image_data[143]), .Y(n5304) );
  AOI22XL U5994 ( .A0(n5558), .A1(image_data[23]), .B0(n5557), .B1(
        image_data[151]), .Y(n5300) );
  AOI22XL U5995 ( .A0(n5546), .A1(image_data[7]), .B0(n5545), .B1(
        image_data[135]), .Y(n5296) );
  AOI22XL U5996 ( .A0(n5582), .A1(image_data[287]), .B0(n5581), .B1(
        image_data[415]), .Y(n5288) );
  AOI22XL U5997 ( .A0(n5570), .A1(image_data[271]), .B0(n5569), .B1(
        image_data[399]), .Y(n5284) );
  AOI22XL U5998 ( .A0(n5558), .A1(image_data[279]), .B0(n5557), .B1(
        image_data[407]), .Y(n5280) );
  NAND2BXL U5999 ( .AN(cmd_reg[1]), .B(n8531), .Y(n6311) );
  NAND2XL U6000 ( .A(cmd_reg[0]), .B(cmd_reg[1]), .Y(n6310) );
  INVXL U6001 ( .A(n7041), .Y(n6620) );
  NOR2XL U6002 ( .A(op4[4]), .B(op4[5]), .Y(n6353) );
  AOI22XL U6003 ( .A0(n7032), .A1(n7040), .B0(n3398), .B1(n7020), .Y(n7023) );
  NAND4XL U6004 ( .A(n8419), .B(n7620), .C(n8393), .D(n8184), .Y(n7020) );
  NAND3XL U6005 ( .A(n8393), .B(n3399), .C(n8184), .Y(n6175) );
  NOR3XL U6006 ( .A(n3379), .B(n8512), .C(n8259), .Y(n4592) );
  NOR3XL U6007 ( .A(n8398), .B(n3379), .C(n8404), .Y(n7097) );
  AOI22XL U6008 ( .A0(n3438), .A1(n6777), .B0(n6767), .B1(n6766), .Y(n6704) );
  INVX1 U6009 ( .A(n5929), .Y(n6767) );
  NAND2XL U6010 ( .A(n7620), .B(n8454), .Y(n7014) );
  AOI22XL U6011 ( .A0(n7096), .A1(n3410), .B0(n3398), .B1(n6768), .Y(n6770) );
  AOI211XL U6012 ( .A0(n6767), .A1(n6766), .B0(n8530), .C0(n8528), .Y(n6768)
         );
  NOR3XL U6013 ( .A(n8452), .B(n8200), .C(n3382), .Y(n5709) );
  NAND2XL U6014 ( .A(n6646), .B(n6984), .Y(n6616) );
  NAND2XL U6015 ( .A(n5921), .B(n6627), .Y(n6625) );
  INVXL U6016 ( .A(n6721), .Y(n5921) );
  NAND2XL U6017 ( .A(n6281), .B(n6984), .Y(n6627) );
  AOI22XL U6018 ( .A0(n6986), .A1(n7008), .B0(n3398), .B1(n6720), .Y(n6723) );
  AOI21XL U6019 ( .A0(n6986), .A1(n6779), .B0(n6778), .Y(n6782) );
  AOI211XL U6020 ( .A0(n3438), .A1(n6777), .B0(n3363), .C0(n6776), .Y(n6778)
         );
  INVXL U6021 ( .A(n6984), .Y(n6776) );
  AND3XL U6022 ( .A(n8529), .B(op2[1]), .C(op2[2]), .Y(n3400) );
  INVXL U6023 ( .A(n6710), .Y(n6639) );
  NAND3XL U6024 ( .A(n8275), .B(n8202), .C(n6341), .Y(n6689) );
  AOI2BB1XL U6025 ( .A0N(n6689), .A1N(n7898), .B0(n3363), .Y(n6687) );
  AOI21XL U6026 ( .A0(n7034), .A1(n6748), .B0(n6776), .Y(n6338) );
  NOR3XL U6027 ( .A(n3377), .B(n6143), .C(n3383), .Y(n6160) );
  INVXL U6028 ( .A(n5698), .Y(n5604) );
  NOR3XL U6029 ( .A(op2[1]), .B(n8528), .C(n6776), .Y(n6720) );
  AOI22XL U6030 ( .A0(n3438), .A1(n6777), .B0(n6728), .B1(n6710), .Y(n6711) );
  AOI22XL U6031 ( .A0(n3410), .A1(n6760), .B0(n3398), .B1(n6638), .Y(n6643) );
  AOI211XL U6032 ( .A0(n6728), .A1(n6710), .B0(n8530), .C0(n8528), .Y(n6638)
         );
  AOI21XL U6033 ( .A0(n7040), .A1(n6760), .B0(n6759), .Y(n6763) );
  AOI31XL U6034 ( .A0(n6758), .A1(n8130), .A2(n3397), .B0(n3363), .Y(n6759) );
  NAND2XL U6035 ( .A(n8467), .B(n6991), .Y(n6758) );
  AOI31XL U6036 ( .A0(n8349), .A1(n8351), .A2(n6758), .B0(n3363), .Y(n6343) );
  AOI21XL U6037 ( .A0(n6994), .A1(n6871), .B0(n6749), .Y(n6752) );
  AOI211XL U6038 ( .A0(n7034), .A1(n6748), .B0(n3363), .C0(n6747), .Y(n6749)
         );
  INVXL U6039 ( .A(n6786), .Y(n6374) );
  AOI21XL U6040 ( .A0(n6994), .A1(n7031), .B0(n6375), .Y(n6785) );
  AOI21XL U6041 ( .A0(n8500), .A1(n6374), .B0(n3363), .Y(n6375) );
  NAND2X1 U6042 ( .A(n6699), .B(n6991), .Y(n6634) );
  INVXL U6043 ( .A(n6389), .Y(n6631) );
  NOR2XL U6044 ( .A(n3438), .B(n6728), .Y(n6391) );
  INVX1 U6045 ( .A(n6747), .Y(n6991) );
  NOR3XL U6046 ( .A(n3431), .B(n3380), .C(n8238), .Y(n6167) );
  NAND3XL U6047 ( .A(n7925), .B(n8349), .C(n8310), .Y(n6735) );
  NOR3XL U6048 ( .A(n3381), .B(n5908), .C(n8228), .Y(n5910) );
  NOR2XL U6049 ( .A(n6777), .B(n6747), .Y(n6389) );
  NAND3XL U6050 ( .A(n8136), .B(n8282), .C(n8317), .Y(n5607) );
  NOR2XL U6051 ( .A(n3438), .B(n6726), .Y(n5700) );
  NAND3XL U6052 ( .A(n8317), .B(n8023), .C(n8125), .Y(n5916) );
  AOI21XL U6053 ( .A0(n7040), .A1(n6734), .B0(n6349), .Y(n6673) );
  AOI31XL U6054 ( .A0(n8023), .A1(n8381), .A2(n6348), .B0(n3363), .Y(n6349) );
  NOR2XL U6055 ( .A(n6401), .B(n5009), .Y(n6151) );
  INVX1 U6056 ( .A(n6902), .Y(n6647) );
  NAND2XL U6057 ( .A(n8467), .B(n6647), .Y(n6348) );
  NAND2XL U6058 ( .A(n6647), .B(n6646), .Y(n6658) );
  INVXL U6059 ( .A(n6791), .Y(n6697) );
  ADDFX2 U6060 ( .A(DP_OP_2677J1_122_9848_n18), .B(DP_OP_2677J1_122_9848_n20), 
        .CI(n6261), .CO(n5897), .S(n6262) );
  NOR4XL U6061 ( .A(n6216), .B(n6215), .C(n6214), .D(n6213), .Y(n6217) );
  NAND4XL U6062 ( .A(n6204), .B(n6203), .C(n6202), .D(n6201), .Y(n6215) );
  NAND4XL U6063 ( .A(n6200), .B(n6199), .C(n6198), .D(n6197), .Y(n6216) );
  NAND4XL U6064 ( .A(n6212), .B(n6211), .C(n6210), .D(n6209), .Y(n6213) );
  NOR4XL U6065 ( .A(n6196), .B(n6195), .C(n6194), .D(n6193), .Y(n6218) );
  NAND4XL U6066 ( .A(n6180), .B(n6179), .C(n6178), .D(n6177), .Y(n6196) );
  NAND4XL U6067 ( .A(n6184), .B(n6183), .C(n6182), .D(n6181), .Y(n6195) );
  NAND4XL U6068 ( .A(n6192), .B(n6191), .C(n6190), .D(n6189), .Y(n6193) );
  AOI22XL U6069 ( .A0(n6574), .A1(n6260), .B0(n6259), .B1(n6571), .Y(n6263) );
  NOR4XL U6070 ( .A(n6238), .B(n6237), .C(n6236), .D(n6235), .Y(n6260) );
  NOR4XL U6071 ( .A(n6258), .B(n6257), .C(n6256), .D(n6255), .Y(n6259) );
  NAND4XL U6072 ( .A(n6226), .B(n6225), .C(n6224), .D(n6223), .Y(n6237) );
  INVXL U6073 ( .A(n5914), .Y(n6030) );
  NAND2XL U6074 ( .A(n6647), .B(n6281), .Y(n6655) );
  NAND2BXL U6075 ( .AN(n6792), .B(n6697), .Y(n6698) );
  NOR2XL U6076 ( .A(n6777), .B(n6902), .Y(n6792) );
  INVXL U6077 ( .A(n6777), .Y(n6780) );
  NAND2XL U6078 ( .A(n8524), .B(n6647), .Y(n5914) );
  AOI22XL U6079 ( .A0(n6574), .A1(n6573), .B0(n6572), .B1(n6571), .Y(n6578) );
  NOR4XL U6080 ( .A(n6518), .B(n6517), .C(n6516), .D(n6515), .Y(n6573) );
  NOR4XL U6081 ( .A(n6570), .B(n6569), .C(n6568), .D(n6567), .Y(n6572) );
  NAND4XL U6082 ( .A(n6502), .B(n6501), .C(n6500), .D(n6499), .Y(n6518) );
  AOI22XL U6083 ( .A0(N2760), .A1(n6418), .B0(N2784), .B1(n6417), .Y(n5269) );
  NOR3XL U6084 ( .A(n8529), .B(op2[1]), .C(op2[2]), .Y(n6750) );
  NAND4XL U6085 ( .A(n8059), .B(n3405), .C(n8370), .D(n8217), .Y(n6870) );
  NOR4XL U6086 ( .A(n5080), .B(n5079), .C(n5078), .D(n5077), .Y(n5081) );
  NAND4XL U6087 ( .A(n5068), .B(n5067), .C(n5066), .D(n5065), .Y(n5079) );
  NAND4XL U6088 ( .A(n5064), .B(n5063), .C(n5062), .D(n5061), .Y(n5080) );
  NAND4XL U6089 ( .A(n5076), .B(n5075), .C(n5074), .D(n5073), .Y(n5077) );
  NOR4XL U6090 ( .A(n5060), .B(n5059), .C(n5058), .D(n5057), .Y(n5082) );
  NAND4XL U6091 ( .A(n5035), .B(n5034), .C(n5033), .D(n5032), .Y(n5059) );
  NAND4XL U6092 ( .A(n5029), .B(n5028), .C(n5027), .D(n5026), .Y(n5060) );
  NAND4XL U6093 ( .A(n5056), .B(n5055), .C(n5054), .D(n5053), .Y(n5057) );
  AOI22XL U6094 ( .A0(n5015), .A1(n3465), .B0(n5014), .B1(n3450), .Y(n5000) );
  AOI22XL U6095 ( .A0(n5012), .A1(n5165), .B0(n5011), .B1(op4[5]), .Y(n5001)
         );
  AOI22XL U6096 ( .A0(n6574), .A1(n5254), .B0(n5253), .B1(n6571), .Y(n5264) );
  NOR4XL U6097 ( .A(n5232), .B(n5231), .C(n5230), .D(n5229), .Y(n5254) );
  NOR4XL U6098 ( .A(n5252), .B(n5251), .C(n5250), .D(n5249), .Y(n5253) );
  NAND4XL U6099 ( .A(n5207), .B(n5206), .C(n5205), .D(n5204), .Y(n5231) );
  NOR4XL U6100 ( .A(n3841), .B(n3840), .C(n3839), .D(n3838), .Y(n3863) );
  NOR4XL U6101 ( .A(n3861), .B(n3860), .C(n3859), .D(n3858), .Y(n3862) );
  NAND4XL U6102 ( .A(n3829), .B(n3828), .C(n3827), .D(n3826), .Y(n3840) );
  CLKINVX2 U6103 ( .A(n7034), .Y(n6646) );
  NAND4XL U6104 ( .A(n4458), .B(n4457), .C(n4456), .D(n4455), .Y(n4469) );
  NOR4XL U6105 ( .A(n3663), .B(n3662), .C(n3661), .D(n3660), .Y(n3685) );
  NOR4XL U6106 ( .A(n3683), .B(n3682), .C(n3681), .D(n3680), .Y(n3684) );
  NAND4XL U6107 ( .A(n3659), .B(n3658), .C(n3657), .D(n3656), .Y(n3660) );
  AOI22XL U6108 ( .A0(n6802), .A1(n6801), .B0(n6800), .B1(n7029), .Y(n6803) );
  AOI22XL U6109 ( .A0(n6574), .A1(n6014), .B0(n6013), .B1(n6571), .Y(n6017) );
  NOR4XL U6110 ( .A(n5992), .B(n5991), .C(n5990), .D(n5989), .Y(n6014) );
  NOR4XL U6111 ( .A(n6012), .B(n6011), .C(n6010), .D(n6009), .Y(n6013) );
  NAND4XL U6112 ( .A(n5988), .B(n5987), .C(n5986), .D(n5985), .Y(n5989) );
  AOI22XL U6113 ( .A0(n6498), .A1(n5972), .B0(n5971), .B1(n6495), .Y(n6018) );
  NOR4XL U6114 ( .A(n5950), .B(n5949), .C(n5948), .D(n5947), .Y(n5972) );
  NOR4XL U6115 ( .A(n5970), .B(n5969), .C(n5968), .D(n5967), .Y(n5971) );
  NAND4XL U6116 ( .A(n5946), .B(n5945), .C(n5944), .D(n5943), .Y(n5947) );
  ADDFX2 U6117 ( .A(DP_OP_2677J1_122_9848_n12), .B(DP_OP_2677J1_122_9848_n14), 
        .CI(n6015), .CO(n6575), .S(n6016) );
  AOI22X1 U6118 ( .A0(n3450), .A1(n4450), .B0(n4449), .B1(n4959), .Y(N2756) );
  NOR4XL U6119 ( .A(n4421), .B(n4420), .C(n4419), .D(n4418), .Y(n4450) );
  NOR4XL U6120 ( .A(n4448), .B(n4447), .C(n4446), .D(n4445), .Y(n4449) );
  NAND4XL U6121 ( .A(n4409), .B(n4408), .C(n4407), .D(n4406), .Y(n4420) );
  AOI22X2 U6122 ( .A0(n5165), .A1(n4064), .B0(n4063), .B1(n4777), .Y(N2780) );
  NAND4XL U6123 ( .A(n4026), .B(n4025), .C(n4024), .D(n4023), .Y(n4042) );
  CLKINVX2 U6124 ( .A(n6800), .Y(n6699) );
  NOR2XL U6125 ( .A(n3376), .B(n8032), .Y(n7010) );
  AOI221XL U6126 ( .A0(n6416), .A1(n6029), .B0(n6415), .B1(n6028), .C0(n6027), 
        .Y(n6346) );
  NAND4XL U6127 ( .A(n4283), .B(n4282), .C(n4281), .D(n4280), .Y(n4294) );
  BUFX1 U6128 ( .A(n4107), .Y(n8568) );
  AOI22XL U6129 ( .A0(op4[5]), .A1(n4106), .B0(n4105), .B1(n8525), .Y(n4107)
         );
  NOR4XL U6130 ( .A(n4084), .B(n4083), .C(n4082), .D(n4081), .Y(n4106) );
  NOR4XL U6131 ( .A(n4104), .B(n4103), .C(n4102), .D(n4101), .Y(n4105) );
  INVX1 U6132 ( .A(N2756), .Y(n5806) );
  NOR4XL U6133 ( .A(n4805), .B(n4804), .C(n4803), .D(n4802), .Y(n4827) );
  NOR4XL U6134 ( .A(n4825), .B(n4824), .C(n4823), .D(n4822), .Y(n4826) );
  NAND4XL U6135 ( .A(n4789), .B(n4788), .C(n4787), .D(n4786), .Y(n4805) );
  NOR4XL U6136 ( .A(n4615), .B(n4614), .C(n4613), .D(n4612), .Y(n4637) );
  NAND4XL U6137 ( .A(n4203), .B(n4202), .C(n4201), .D(n4200), .Y(n4209) );
  NAND4XL U6138 ( .A(n3988), .B(n3987), .C(n3986), .D(n3985), .Y(n3999) );
  NOR4XL U6139 ( .A(n4337), .B(n4336), .C(n4335), .D(n4334), .Y(n4359) );
  NOR4XL U6140 ( .A(n4357), .B(n4356), .C(n4355), .D(n4354), .Y(n4358) );
  NAND4XL U6141 ( .A(n4321), .B(n4320), .C(n4319), .D(n4318), .Y(n4337) );
  AOI22XL U6142 ( .A0(op4[5]), .A1(n3727), .B0(n3726), .B1(n8525), .Y(n3728)
         );
  NOR4XL U6143 ( .A(n3705), .B(n3704), .C(n3703), .D(n3702), .Y(n3727) );
  NOR4XL U6144 ( .A(n3725), .B(n3724), .C(n3723), .D(n3722), .Y(n3726) );
  NAND2XL U6145 ( .A(n8432), .B(n8419), .Y(n7016) );
  NAND2XL U6146 ( .A(n6819), .B(op4[3]), .Y(n6824) );
  NAND4XL U6147 ( .A(n3873), .B(n3872), .C(n3871), .D(n3870), .Y(n3905) );
  BUFX1 U6148 ( .A(n3980), .Y(n8569) );
  AOI22XL U6149 ( .A0(op4[5]), .A1(n3979), .B0(n3978), .B1(n8525), .Y(n3980)
         );
  NOR4XL U6150 ( .A(n3957), .B(n3956), .C(n3955), .D(n3954), .Y(n3979) );
  NOR4XL U6151 ( .A(n3977), .B(n3976), .C(n3975), .D(n3974), .Y(n3978) );
  AOI22XL U6152 ( .A0(N2759), .A1(n6418), .B0(N2783), .B1(n6417), .Y(n6176) );
  INVXL U6153 ( .A(N2758), .Y(n5705) );
  NAND4XL U6154 ( .A(n4363), .B(n4362), .C(n4361), .D(n4360), .Y(n4379) );
  NOR2XL U6155 ( .A(n8531), .B(n6027), .Y(n4593) );
  NOR2XL U6156 ( .A(cmd_reg[0]), .B(n6027), .Y(n4594) );
  AOI31XL U6157 ( .A0(n7041), .A1(n8419), .A2(n8440), .B0(n3363), .Y(n7042) );
  NOR2XL U6158 ( .A(cmd_reg[3]), .B(n6583), .Y(n6313) );
  INVXL U6159 ( .A(n6383), .Y(n6299) );
  AOI22XL U6160 ( .A0(n5546), .A1(image_data[256]), .B0(n5545), .B1(
        image_data[384]), .Y(n5486) );
  AOI22XL U6161 ( .A0(n5552), .A1(image_data[352]), .B0(n5551), .B1(
        image_data[480]), .Y(n5483) );
  AOI22XL U6162 ( .A0(n5548), .A1(image_data[320]), .B0(n5547), .B1(
        image_data[448]), .Y(n5485) );
  AOI22XL U6163 ( .A0(n5550), .A1(image_data[288]), .B0(n5549), .B1(
        image_data[416]), .Y(n5484) );
  NAND4XL U6164 ( .A(n5506), .B(n5505), .C(n5504), .D(n5503), .Y(n5522) );
  AOI22XL U6165 ( .A0(n5550), .A1(image_data[32]), .B0(n5549), .B1(
        image_data[160]), .Y(n5504) );
  AOI22XL U6166 ( .A0(n5548), .A1(image_data[64]), .B0(n5547), .B1(
        image_data[192]), .Y(n5505) );
  AOI22XL U6167 ( .A0(n5552), .A1(image_data[96]), .B0(n5551), .B1(
        image_data[224]), .Y(n5503) );
  NAND4XL U6168 ( .A(n5490), .B(n5489), .C(n5488), .D(n5487), .Y(n5501) );
  AOI22XL U6169 ( .A0(n5560), .A1(image_data[336]), .B0(n5559), .B1(
        image_data[464]), .Y(n5489) );
  AOI22XL U6170 ( .A0(n5562), .A1(image_data[304]), .B0(n5561), .B1(
        image_data[432]), .Y(n5488) );
  AOI22XL U6171 ( .A0(n5564), .A1(image_data[368]), .B0(n5563), .B1(
        image_data[496]), .Y(n5487) );
  AOI22XL U6172 ( .A0(n5546), .A1(image_data[257]), .B0(n5545), .B1(
        image_data[385]), .Y(n5402) );
  AOI22XL U6173 ( .A0(n5552), .A1(image_data[353]), .B0(n5551), .B1(
        image_data[481]), .Y(n5399) );
  AOI22XL U6174 ( .A0(n5548), .A1(image_data[321]), .B0(n5547), .B1(
        image_data[449]), .Y(n5401) );
  AOI22XL U6175 ( .A0(n5550), .A1(image_data[289]), .B0(n5549), .B1(
        image_data[417]), .Y(n5400) );
  NAND4XL U6176 ( .A(n5422), .B(n5421), .C(n5420), .D(n5419), .Y(n5438) );
  AOI22XL U6177 ( .A0(n5550), .A1(image_data[33]), .B0(n5549), .B1(
        image_data[161]), .Y(n5420) );
  AOI22XL U6178 ( .A0(n5548), .A1(image_data[65]), .B0(n5547), .B1(
        image_data[193]), .Y(n5421) );
  AOI22XL U6179 ( .A0(n5552), .A1(image_data[97]), .B0(n5551), .B1(
        image_data[225]), .Y(n5419) );
  NAND4XL U6180 ( .A(n5406), .B(n5405), .C(n5404), .D(n5403), .Y(n5417) );
  AOI22XL U6181 ( .A0(n5560), .A1(image_data[337]), .B0(n5559), .B1(
        image_data[465]), .Y(n5405) );
  AOI22XL U6182 ( .A0(n5562), .A1(image_data[305]), .B0(n5561), .B1(
        image_data[433]), .Y(n5404) );
  AOI22XL U6183 ( .A0(n5564), .A1(image_data[369]), .B0(n5563), .B1(
        image_data[497]), .Y(n5403) );
  AOI22XL U6184 ( .A0(n5546), .A1(image_data[258]), .B0(n5545), .B1(
        image_data[386]), .Y(n4540) );
  AOI22XL U6185 ( .A0(n5552), .A1(image_data[354]), .B0(n5551), .B1(
        image_data[482]), .Y(n4537) );
  AOI22XL U6186 ( .A0(n5548), .A1(image_data[322]), .B0(n5547), .B1(
        image_data[450]), .Y(n4539) );
  AOI22XL U6187 ( .A0(n5550), .A1(image_data[290]), .B0(n5549), .B1(
        image_data[418]), .Y(n4538) );
  NAND4XL U6188 ( .A(n4568), .B(n4567), .C(n4566), .D(n4565), .Y(n4584) );
  AOI22XL U6189 ( .A0(n5550), .A1(image_data[34]), .B0(n5549), .B1(
        image_data[162]), .Y(n4566) );
  AOI22XL U6190 ( .A0(n5548), .A1(image_data[66]), .B0(n5547), .B1(
        image_data[194]), .Y(n4567) );
  AOI22XL U6191 ( .A0(n5552), .A1(image_data[98]), .B0(n5551), .B1(
        image_data[226]), .Y(n4565) );
  NAND4XL U6192 ( .A(n4544), .B(n4543), .C(n4542), .D(n4541), .Y(n4563) );
  AOI22XL U6193 ( .A0(n5560), .A1(image_data[338]), .B0(n5559), .B1(
        image_data[466]), .Y(n4543) );
  AOI22XL U6194 ( .A0(n5562), .A1(image_data[306]), .B0(n5561), .B1(
        image_data[434]), .Y(n4542) );
  AOI22XL U6195 ( .A0(n5564), .A1(image_data[370]), .B0(n5563), .B1(
        image_data[498]), .Y(n4541) );
  AOI22XL U6196 ( .A0(n5546), .A1(image_data[259]), .B0(n5545), .B1(
        image_data[387]), .Y(n5528) );
  AOI22XL U6197 ( .A0(n5552), .A1(image_data[355]), .B0(n5551), .B1(
        image_data[483]), .Y(n5525) );
  AOI22XL U6198 ( .A0(n5548), .A1(image_data[323]), .B0(n5547), .B1(
        image_data[451]), .Y(n5527) );
  AOI22XL U6199 ( .A0(n5550), .A1(image_data[291]), .B0(n5549), .B1(
        image_data[419]), .Y(n5526) );
  NAND4XL U6200 ( .A(n5556), .B(n5555), .C(n5554), .D(n5553), .Y(n5596) );
  AOI22XL U6201 ( .A0(n5550), .A1(image_data[35]), .B0(n5549), .B1(
        image_data[163]), .Y(n5554) );
  AOI22XL U6202 ( .A0(n5548), .A1(image_data[67]), .B0(n5547), .B1(
        image_data[195]), .Y(n5555) );
  AOI22XL U6203 ( .A0(n5552), .A1(image_data[99]), .B0(n5551), .B1(
        image_data[227]), .Y(n5553) );
  NAND4XL U6204 ( .A(n5532), .B(n5531), .C(n5530), .D(n5529), .Y(n5543) );
  AOI22XL U6205 ( .A0(n5560), .A1(image_data[339]), .B0(n5559), .B1(
        image_data[467]), .Y(n5531) );
  AOI22XL U6206 ( .A0(n5562), .A1(image_data[307]), .B0(n5561), .B1(
        image_data[435]), .Y(n5530) );
  AOI22XL U6207 ( .A0(n5564), .A1(image_data[371]), .B0(n5563), .B1(
        image_data[499]), .Y(n5529) );
  AOI22XL U6208 ( .A0(n5546), .A1(image_data[260]), .B0(n5545), .B1(
        image_data[388]), .Y(n5444) );
  AOI22XL U6209 ( .A0(n5552), .A1(image_data[356]), .B0(n5551), .B1(
        image_data[484]), .Y(n5441) );
  AOI22XL U6210 ( .A0(n5548), .A1(image_data[324]), .B0(n5547), .B1(
        image_data[452]), .Y(n5443) );
  AOI22XL U6211 ( .A0(n5550), .A1(image_data[292]), .B0(n5549), .B1(
        image_data[420]), .Y(n5442) );
  NAND4XL U6212 ( .A(n5464), .B(n5463), .C(n5462), .D(n5461), .Y(n5480) );
  AOI22XL U6213 ( .A0(n5550), .A1(image_data[36]), .B0(n5549), .B1(
        image_data[164]), .Y(n5462) );
  AOI22XL U6214 ( .A0(n5548), .A1(image_data[68]), .B0(n5547), .B1(
        image_data[196]), .Y(n5463) );
  AOI22XL U6215 ( .A0(n5552), .A1(image_data[100]), .B0(n5551), .B1(
        image_data[228]), .Y(n5461) );
  NAND4XL U6216 ( .A(n5448), .B(n5447), .C(n5446), .D(n5445), .Y(n5459) );
  AOI22XL U6217 ( .A0(n5560), .A1(image_data[340]), .B0(n5559), .B1(
        image_data[468]), .Y(n5447) );
  AOI22XL U6218 ( .A0(n5562), .A1(image_data[308]), .B0(n5561), .B1(
        image_data[436]), .Y(n5446) );
  AOI22XL U6219 ( .A0(n5564), .A1(image_data[372]), .B0(n5563), .B1(
        image_data[500]), .Y(n5445) );
  AOI22XL U6220 ( .A0(n5546), .A1(image_data[261]), .B0(n5545), .B1(
        image_data[389]), .Y(n5360) );
  AOI22XL U6221 ( .A0(n5552), .A1(image_data[357]), .B0(n5551), .B1(
        image_data[485]), .Y(n5357) );
  AOI22XL U6222 ( .A0(n5548), .A1(image_data[325]), .B0(n5547), .B1(
        image_data[453]), .Y(n5359) );
  AOI22XL U6223 ( .A0(n5550), .A1(image_data[293]), .B0(n5549), .B1(
        image_data[421]), .Y(n5358) );
  NAND4XL U6224 ( .A(n5380), .B(n5379), .C(n5378), .D(n5377), .Y(n5396) );
  AOI22XL U6225 ( .A0(n5550), .A1(image_data[37]), .B0(n5549), .B1(
        image_data[165]), .Y(n5378) );
  AOI22XL U6226 ( .A0(n5548), .A1(image_data[69]), .B0(n5547), .B1(
        image_data[197]), .Y(n5379) );
  AOI22XL U6227 ( .A0(n5552), .A1(image_data[101]), .B0(n5551), .B1(
        image_data[229]), .Y(n5377) );
  NAND4XL U6228 ( .A(n5364), .B(n5363), .C(n5362), .D(n5361), .Y(n5375) );
  AOI22XL U6229 ( .A0(n5560), .A1(image_data[341]), .B0(n5559), .B1(
        image_data[469]), .Y(n5363) );
  AOI22XL U6230 ( .A0(n5562), .A1(image_data[309]), .B0(n5561), .B1(
        image_data[437]), .Y(n5362) );
  AOI22XL U6231 ( .A0(n5564), .A1(image_data[373]), .B0(n5563), .B1(
        image_data[501]), .Y(n5361) );
  AOI22XL U6232 ( .A0(n5546), .A1(image_data[262]), .B0(n5545), .B1(
        image_data[390]), .Y(n5318) );
  AOI22XL U6233 ( .A0(n5552), .A1(image_data[358]), .B0(n5551), .B1(
        image_data[486]), .Y(n5315) );
  AOI22XL U6234 ( .A0(n5548), .A1(image_data[326]), .B0(n5547), .B1(
        image_data[454]), .Y(n5317) );
  AOI22XL U6235 ( .A0(n5550), .A1(image_data[294]), .B0(n5549), .B1(
        image_data[422]), .Y(n5316) );
  NAND4XL U6236 ( .A(n5338), .B(n5337), .C(n5336), .D(n5335), .Y(n5354) );
  AOI22XL U6237 ( .A0(n5550), .A1(image_data[38]), .B0(n5549), .B1(
        image_data[166]), .Y(n5336) );
  AOI22XL U6238 ( .A0(n5548), .A1(image_data[70]), .B0(n5547), .B1(
        image_data[198]), .Y(n5337) );
  AOI22XL U6239 ( .A0(n5552), .A1(image_data[102]), .B0(n5551), .B1(
        image_data[230]), .Y(n5335) );
  NAND4XL U6240 ( .A(n5322), .B(n5321), .C(n5320), .D(n5319), .Y(n5333) );
  AOI22XL U6241 ( .A0(n5560), .A1(image_data[342]), .B0(n5559), .B1(
        image_data[470]), .Y(n5321) );
  AOI22XL U6242 ( .A0(n5562), .A1(image_data[310]), .B0(n5561), .B1(
        image_data[438]), .Y(n5320) );
  AOI22XL U6243 ( .A0(n5564), .A1(image_data[374]), .B0(n5563), .B1(
        image_data[502]), .Y(n5319) );
  AOI22XL U6244 ( .A0(n5546), .A1(image_data[263]), .B0(n5545), .B1(
        image_data[391]), .Y(n5276) );
  AOI22XL U6245 ( .A0(n5552), .A1(image_data[359]), .B0(n5551), .B1(
        image_data[487]), .Y(n5273) );
  AOI22XL U6246 ( .A0(n5548), .A1(image_data[327]), .B0(n5547), .B1(
        image_data[455]), .Y(n5275) );
  AOI22XL U6247 ( .A0(n5550), .A1(image_data[295]), .B0(n5549), .B1(
        image_data[423]), .Y(n5274) );
  NAND4XL U6248 ( .A(n5296), .B(n5295), .C(n5294), .D(n5293), .Y(n5312) );
  AOI22XL U6249 ( .A0(n5550), .A1(image_data[39]), .B0(n5549), .B1(
        image_data[167]), .Y(n5294) );
  AOI22XL U6250 ( .A0(n5548), .A1(image_data[71]), .B0(n5547), .B1(
        image_data[199]), .Y(n5295) );
  AOI22XL U6251 ( .A0(n5552), .A1(image_data[103]), .B0(n5551), .B1(
        image_data[231]), .Y(n5293) );
  NAND4XL U6252 ( .A(n5280), .B(n5279), .C(n5278), .D(n5277), .Y(n5291) );
  AOI22XL U6253 ( .A0(n5560), .A1(image_data[343]), .B0(n5559), .B1(
        image_data[471]), .Y(n5279) );
  AOI22XL U6254 ( .A0(n5562), .A1(image_data[311]), .B0(n5561), .B1(
        image_data[439]), .Y(n5278) );
  AOI22XL U6255 ( .A0(n5564), .A1(image_data[375]), .B0(n5563), .B1(
        image_data[503]), .Y(n5277) );
  INVXL U6256 ( .A(n4588), .Y(n8468) );
  NOR2X1 U6257 ( .A(cmd_reg[2]), .B(n6310), .Y(n8466) );
  INVXL U6258 ( .A(n6313), .Y(n6312) );
  NAND2XL U6259 ( .A(IROM_A[3]), .B(n8487), .Y(n8486) );
  INVXL U6260 ( .A(n8477), .Y(n8465) );
  OAI22XL U6261 ( .A0(in_done), .A1(n8523), .B0(n8489), .B1(n8534), .Y(n8478)
         );
  NAND2XL U6262 ( .A(IROM_A[0]), .B(n8478), .Y(n8477) );
  NOR2XL U6263 ( .A(n6299), .B(op4[3]), .Y(n6386) );
  NOR3XL U6264 ( .A(n6312), .B(cmd_reg[2]), .C(n6415), .Y(n6383) );
  NAND2XL U6265 ( .A(IROM_A[1]), .B(n8465), .Y(n8464) );
  NOR2XL U6266 ( .A(n8519), .B(n8464), .Y(n8487) );
  NOR2XL U6267 ( .A(n8527), .B(n8486), .Y(n6382) );
  INVXL U6268 ( .A(n6382), .Y(n8479) );
  NOR2XL U6269 ( .A(done), .B(n8489), .Y(n6322) );
  NOR2XL U6270 ( .A(n8481), .B(n8489), .Y(n8488) );
  NAND2BXL U6271 ( .AN(in_done), .B(n8480), .Y(n8463) );
  AOI21XL U6272 ( .A0(n7032), .A1(n6688), .B0(n6621), .Y(n8084) );
  AOI21XL U6273 ( .A0(n8080), .A1(n3399), .B0(n3363), .Y(n6621) );
  NOR2XL U6274 ( .A(n6620), .B(n8182), .Y(n8080) );
  NOR2BX1 U6275 ( .AN(n8080), .B(n8084), .Y(n8188) );
  NOR3XL U6276 ( .A(n8513), .B(n8182), .C(n8368), .Y(n6970) );
  INVXL U6277 ( .A(n8371), .Y(n8099) );
  AOI21XL U6278 ( .A0(n6970), .A1(n8101), .B0(n3363), .Y(n5930) );
  NAND2XL U6279 ( .A(n6970), .B(n8096), .Y(n8371) );
  AOI211XL U6280 ( .A0(n7029), .A1(n7034), .B0(n3363), .C0(n7033), .Y(n7030)
         );
  CLKINVX2 U6281 ( .A(n3417), .Y(n8413) );
  NOR2X2 U6282 ( .A(n6802), .B(n7029), .Y(n8511) );
  AOI2BB1XL U6283 ( .A0N(n5811), .A1N(n8398), .B0(n3363), .Y(n5810) );
  AOI21XL U6284 ( .A0(n7032), .A1(n7008), .B0(n7007), .Y(n7009) );
  AOI31XL U6285 ( .A0(n7010), .A1(n7995), .A2(n8406), .B0(n3363), .Y(n7007) );
  INVXL U6286 ( .A(n7750), .Y(n8089) );
  CLKINVX2 U6287 ( .A(n6978), .Y(n8086) );
  AOI21XL U6288 ( .A0(n6975), .A1(n8454), .B0(n3363), .Y(n6356) );
  NAND2XL U6289 ( .A(n6975), .B(n8086), .Y(n7750) );
  AOI2BB1XL U6290 ( .A0N(n7016), .A1N(n7014), .B0(n3363), .Y(n7015) );
  CLKINVX2 U6291 ( .A(n7747), .Y(n8433) );
  CLKINVX2 U6292 ( .A(n7023), .Y(n8420) );
  INVX1 U6293 ( .A(n3407), .Y(n3429) );
  AOI21XL U6294 ( .A0(n7096), .A1(n6688), .B0(n6174), .Y(n6269) );
  AOI2BB1XL U6295 ( .A0N(n6175), .A1N(n8260), .B0(n3363), .Y(n6174) );
  CLKINVX3 U6296 ( .A(n8184), .Y(n8417) );
  CLKINVX2 U6297 ( .A(n6269), .Y(n8091) );
  NAND3XL U6298 ( .A(n8101), .B(n3399), .C(n7684), .Y(n6998) );
  AOI21XL U6299 ( .A0(n7582), .A1(n8425), .B0(n3363), .Y(n6366) );
  INVXL U6300 ( .A(n6998), .Y(n7582) );
  CLKINVX2 U6301 ( .A(n3399), .Y(n8368) );
  CLKINVX2 U6302 ( .A(n8028), .Y(n8018) );
  CLKINVX3 U6303 ( .A(n8101), .Y(n8512) );
  AOI21XL U6304 ( .A0(n4592), .A1(n8209), .B0(n3363), .Y(n4591) );
  CLKINVX2 U6305 ( .A(n7564), .Y(n8426) );
  INVXL U6306 ( .A(n4592), .Y(n7560) );
  INVX1 U6307 ( .A(n7572), .Y(n8410) );
  AOI21XL U6308 ( .A0(n7097), .A1(n8304), .B0(n3363), .Y(n7094) );
  CLKINVX2 U6309 ( .A(n7575), .Y(n8407) );
  NAND2XL U6310 ( .A(n7097), .B(n8407), .Y(n7572) );
  AOI22XL U6311 ( .A0(n8458), .A1(n6418), .B0(n5698), .B1(n6417), .Y(n5699) );
  NAND3XL U6312 ( .A(n7995), .B(n8406), .C(n8304), .Y(n7002) );
  AOI21XL U6313 ( .A0(n7096), .A1(n7008), .B0(n6406), .Y(n7003) );
  AOI2BB1XL U6314 ( .A0N(n7002), .A1N(n8302), .B0(n3363), .Y(n6406) );
  CLKINVX2 U6315 ( .A(n7003), .Y(n7766) );
  CLKINVX2 U6316 ( .A(n6707), .Y(n8388) );
  NAND3XL U6317 ( .A(n7995), .B(n8454), .C(n8387), .Y(n6705) );
  NAND2X1 U6318 ( .A(n6992), .B(n5929), .Y(n7620) );
  BUFX1 U6319 ( .A(n6355), .Y(n8430) );
  NOR2XL U6320 ( .A(n3438), .B(n6767), .Y(n6355) );
  CLKINVX2 U6321 ( .A(n6770), .Y(n8455) );
  INVX1 U6322 ( .A(n3408), .Y(n3428) );
  AOI21XL U6323 ( .A0(n7096), .A1(n7040), .B0(n5708), .Y(n5804) );
  AOI21XL U6324 ( .A0(n5709), .A1(n8202), .B0(n3363), .Y(n5708) );
  CLKINVX3 U6325 ( .A(n7620), .Y(n8452) );
  CLKINVX2 U6326 ( .A(n5804), .Y(n8394) );
  AOI21XL U6327 ( .A0(n6665), .A1(n6668), .B0(n3363), .Y(n6666) );
  INVX1 U6328 ( .A(n8260), .Y(n7684) );
  CLKINVX2 U6329 ( .A(n6683), .Y(n8262) );
  AOI22XL U6330 ( .A0(n6124), .A1(n6418), .B0(n6123), .B1(n6417), .Y(n6125) );
  AOI21XL U6331 ( .A0(n6627), .A1(n6616), .B0(n3363), .Y(n6614) );
  CLKINVX2 U6332 ( .A(n8404), .Y(n8209) );
  AOI22XL U6333 ( .A0(n6986), .A1(n7095), .B0(n3398), .B1(n6625), .Y(n6626) );
  NOR2X1 U6334 ( .A(n6777), .B(n6766), .Y(n8302) );
  CLKINVX3 U6335 ( .A(n8304), .Y(n8207) );
  CLKINVX2 U6336 ( .A(n6723), .Y(n8305) );
  INVX1 U6337 ( .A(n3406), .Y(n3427) );
  CLKINVX2 U6338 ( .A(n6782), .Y(n8364) );
  AOI211XL U6339 ( .A0(n3438), .A1(n8483), .B0(n3363), .C0(n6776), .Y(n6288)
         );
  CLKINVX2 U6340 ( .A(n8287), .Y(n7918) );
  CLKINVX2 U6341 ( .A(n6294), .Y(n7919) );
  AOI21XL U6342 ( .A0(n6986), .A1(n7040), .B0(n6985), .Y(n7569) );
  AOI21XL U6343 ( .A0(n6987), .A1(n6341), .B0(n3363), .Y(n6985) );
  CLKINVX2 U6344 ( .A(n7569), .Y(n8148) );
  NAND2XL U6345 ( .A(n6987), .B(n8148), .Y(n7566) );
  AOI22XL U6346 ( .A0(n6127), .A1(n6420), .B0(n6126), .B1(n6421), .Y(n7445) );
  CLKINVX3 U6347 ( .A(n8202), .Y(n8273) );
  CLKINVX2 U6348 ( .A(n6691), .Y(n8276) );
  AOI21XL U6349 ( .A0(n6760), .A1(n6871), .B0(n6144), .Y(n7987) );
  AOI21XL U6350 ( .A0(n7983), .A1(n8171), .B0(n3363), .Y(n6144) );
  AOI21XL U6351 ( .A0(n6160), .A1(n7907), .B0(n3363), .Y(n6159) );
  CLKINVX2 U6352 ( .A(n6163), .Y(n8172) );
  AOI21XL U6353 ( .A0(n5923), .A1(n7975), .B0(n3363), .Y(n5922) );
  AOI21XL U6354 ( .A0(n6760), .A1(n7008), .B0(n6137), .Y(n7978) );
  AOI21XL U6355 ( .A0(n7972), .A1(n8289), .B0(n3363), .Y(n6137) );
  CLKINVX3 U6356 ( .A(n8177), .Y(n8301) );
  BUFX1 U6357 ( .A(n6138), .Y(n8362) );
  NOR2XL U6358 ( .A(n6777), .B(n6710), .Y(n6138) );
  CLKINVX2 U6359 ( .A(n6714), .Y(n8290) );
  NAND3XL U6360 ( .A(n8289), .B(n8153), .C(n7918), .Y(n6712) );
  AOI22XL U6361 ( .A0(N2774), .A1(n6421), .B0(N2766), .B1(n6420), .Y(n5801) );
  BUFX1 U6362 ( .A(n6289), .Y(n8287) );
  NOR2XL U6363 ( .A(n3438), .B(n6710), .Y(n6289) );
  CLKINVX2 U6364 ( .A(n6643), .Y(n8235) );
  INVX1 U6365 ( .A(n3409), .Y(n3426) );
  CLKINVX2 U6366 ( .A(n6763), .Y(n8358) );
  NOR3X2 U6367 ( .A(n3378), .B(n6763), .C(n6761), .Y(n8361) );
  CLKINVX2 U6368 ( .A(n6678), .Y(n8255) );
  INVXL U6369 ( .A(n6728), .Y(n6142) );
  CLKINVX2 U6370 ( .A(n6143), .Y(n8171) );
  CLKINVX2 U6371 ( .A(n8351), .Y(n7898) );
  CLKINVX2 U6372 ( .A(n6752), .Y(n8352) );
  CLKINVX2 U6373 ( .A(n6785), .Y(n7926) );
  AOI21XL U6374 ( .A0(n6634), .A1(n8500), .B0(n3363), .Y(n6276) );
  NOR2XL U6375 ( .A(n3413), .B(n8499), .Y(n8502) );
  CLKINVX2 U6376 ( .A(n6279), .Y(n8507) );
  CLKINVX2 U6377 ( .A(n8499), .Y(n7975) );
  AOI21XL U6378 ( .A0(n6994), .A1(n7008), .B0(n6632), .Y(n6633) );
  INVX1 U6379 ( .A(n3387), .Y(n8199) );
  NAND2XL U6380 ( .A(n6631), .B(n7878), .Y(n6950) );
  INVXL U6381 ( .A(n6950), .Y(n6964) );
  AOI21XL U6382 ( .A0(n6964), .A1(n8317), .B0(n3363), .Y(n6390) );
  INVXL U6383 ( .A(n6391), .Y(n7878) );
  INVX1 U6384 ( .A(n5700), .Y(n8317) );
  INVXL U6385 ( .A(n3411), .Y(n3412) );
  AOI22XL U6386 ( .A0(n6994), .A1(n3410), .B0(n3398), .B1(n6727), .Y(n7058) );
  AOI22XL U6387 ( .A0(n3438), .A1(n8483), .B0(n6726), .B1(n6728), .Y(n6727) );
  BUFX1 U6388 ( .A(n6391), .Y(n8315) );
  CLKINVX2 U6389 ( .A(n3412), .Y(n8318) );
  NAND3XL U6390 ( .A(n8317), .B(n7878), .C(n8130), .Y(n6729) );
  AOI21XL U6391 ( .A0(n6992), .A1(n6991), .B0(n3380), .Y(n8021) );
  INVXL U6392 ( .A(n7577), .Y(n8134) );
  NAND2XL U6393 ( .A(n8021), .B(n8131), .Y(n7577) );
  AOI21XL U6394 ( .A0(n6688), .A1(n6734), .B0(n6166), .Y(n6170) );
  AOI21XL U6395 ( .A0(n6167), .A1(n8310), .B0(n6337), .Y(n6166) );
  CLKINVX2 U6396 ( .A(n6170), .Y(n8166) );
  AOI2BB1XL U6397 ( .A0N(n6735), .A1N(n8214), .B0(n3363), .Y(n6733) );
  CLKINVX3 U6398 ( .A(n8349), .Y(n3431) );
  CLKINVX2 U6399 ( .A(n7940), .Y(n8311) );
  NOR3XL U6400 ( .A(n5908), .B(n8308), .C(n8214), .Y(n6878) );
  AOI21XL U6401 ( .A0(n6878), .A1(n8159), .B0(n3363), .Y(n6031) );
  CLKINVX3 U6402 ( .A(n7925), .Y(n8308) );
  INVX1 U6403 ( .A(n3433), .Y(n3434) );
  NOR2BXL U6404 ( .AN(n6878), .B(n6884), .Y(n8272) );
  AOI21XL U6405 ( .A0(n7095), .A1(n6734), .B0(n5909), .Y(n7935) );
  NOR3XL U6406 ( .A(n3381), .B(n7888), .C(n3452), .Y(n6592) );
  AOI21XL U6407 ( .A0(n6734), .A1(n7008), .B0(n6324), .Y(n6325) );
  AOI21XL U6408 ( .A0(n6592), .A1(n8282), .B0(n6337), .Y(n6324) );
  CLKINVX2 U6409 ( .A(n6325), .Y(n8137) );
  AOI2BB1XL U6410 ( .A0N(n5607), .A1N(n8490), .B0(n3363), .Y(n5606) );
  AOI21XL U6411 ( .A0(n3410), .A1(n6734), .B0(n5915), .Y(n5919) );
  AOI2BB1XL U6412 ( .A0N(n5916), .A1N(n7513), .B0(n3363), .Y(n5915) );
  BUFX1 U6413 ( .A(n5700), .Y(n7887) );
  CLKINVX2 U6414 ( .A(n5919), .Y(n7698) );
  BUFX1 U6415 ( .A(n8222), .Y(n3455) );
  NOR2XL U6416 ( .A(n6726), .B(n8483), .Y(n8222) );
  CLKINVX2 U6417 ( .A(n6673), .Y(n8224) );
  AOI21XL U6418 ( .A0(n6650), .A1(n6348), .B0(n3363), .Y(n6150) );
  CLKINVX2 U6419 ( .A(n6154), .Y(n8240) );
  AOI21XL U6420 ( .A0(n6904), .A1(n6871), .B0(n6648), .Y(n6649) );
  AND3XL U6421 ( .A(n8267), .B(n6650), .C(n8218), .Y(n8221) );
  AOI22XL U6422 ( .A0(n4871), .A1(n6420), .B0(n8459), .B1(n6421), .Y(n8014) );
  CLKINVX3 U6423 ( .A(n8267), .Y(n8214) );
  AOI21XL U6424 ( .A0(n6655), .A1(n6658), .B0(n3363), .Y(n6656) );
  AOI21XL U6425 ( .A0(n6904), .A1(n7095), .B0(n6282), .Y(n6285) );
  AOI21XL U6426 ( .A0(n6697), .A1(n6655), .B0(n3363), .Y(n6282) );
  NAND2XL U6427 ( .A(n7864), .B(n6655), .Y(n6369) );
  CLKINVX2 U6428 ( .A(n6285), .Y(n7349) );
  NOR2X1 U6429 ( .A(n6285), .B(n6369), .Y(n7352) );
  INVXL U6430 ( .A(n7864), .Y(n8280) );
  CLKINVX2 U6431 ( .A(n6701), .Y(n8283) );
  NOR2XL U6432 ( .A(n6792), .B(n8490), .Y(n8493) );
  CLKINVX2 U6433 ( .A(n6963), .Y(n8498) );
  INVXL U6434 ( .A(n7312), .Y(n8128) );
  NAND2XL U6435 ( .A(n6780), .B(n6825), .Y(n7317) );
  BUFX1 U6436 ( .A(n5605), .Y(n8492) );
  NOR2XL U6437 ( .A(n6777), .B(n5914), .Y(n5605) );
  NAND2XL U6438 ( .A(n8493), .B(n8498), .Y(n7312) );
  AOI22XL U6439 ( .A0(N2757), .A1(n6418), .B0(N2781), .B1(n6417), .Y(n5928) );
  CLKINVX2 U6440 ( .A(n6744), .Y(n8336) );
  AOI2BB1XL U6441 ( .A0N(n6905), .A1N(n8438), .B0(n3363), .Y(n6903) );
  CLKINVX2 U6442 ( .A(n8380), .Y(n7874) );
  CLKINVX3 U6443 ( .A(n6145), .Y(n8111) );
  NOR3XL U6444 ( .A(n8438), .B(n8343), .C(n8378), .Y(n8074) );
  AOI21XL U6445 ( .A0(n8074), .A1(n8370), .B0(n3363), .Y(n6132) );
  CLKINVX3 U6446 ( .A(n8076), .Y(n8378) );
  INVX1 U6447 ( .A(n3435), .Y(n3436) );
  NOR2BXL U6448 ( .AN(n8074), .B(n8079), .Y(n8327) );
  INVXL U6449 ( .A(n7963), .Y(n7261) );
  CLKINVX2 U6450 ( .A(n6875), .Y(n8345) );
  INVXL U6451 ( .A(n8268), .Y(n8376) );
  NAND3XL U6452 ( .A(n8329), .B(n8059), .C(n3405), .Y(n7306) );
  INVXL U6453 ( .A(n7740), .Y(n7690) );
  AOI2BB1XL U6454 ( .A0N(n7306), .A1N(n8511), .B0(n3363), .Y(n5599) );
  CLKINVX3 U6455 ( .A(n8059), .Y(n8513) );
  INVXL U6456 ( .A(n7445), .Y(n7517) );
  INVXL U6457 ( .A(n3421), .Y(n6943) );
  INVXL U6458 ( .A(n7895), .Y(n7902) );
  INVXL U6459 ( .A(n8055), .Y(n7487) );
  NOR2XL U6460 ( .A(n5800), .B(n6583), .Y(n7377) );
  AOI22XL U6461 ( .A0(N2758), .A1(n6418), .B0(N2782), .B1(n6417), .Y(n5800) );
  INVXL U6462 ( .A(n7956), .Y(n7930) );
  INVXL U6463 ( .A(n5812), .Y(n7723) );
  CLKINVX2 U6464 ( .A(n6806), .Y(n8297) );
  NAND3XL U6465 ( .A(n7455), .B(n8412), .C(n8329), .Y(n6804) );
  NOR2X1 U6466 ( .A(n5903), .B(n6583), .Y(n6951) );
  AOI22XL U6467 ( .A0(N2756), .A1(n6418), .B0(N2780), .B1(n6417), .Y(n5903) );
  CLKINVX3 U6468 ( .A(n7455), .Y(n8294) );
  AOI21XL U6469 ( .A0(n7010), .A1(n6795), .B0(n3363), .Y(n6793) );
  AOI21XL U6470 ( .A0(n6400), .A1(n8432), .B0(n3363), .Y(n6399) );
  NAND2XL U6471 ( .A(n6957), .B(n6400), .Y(n8069) );
  CLKINVX2 U6472 ( .A(n5808), .Y(n8509) );
  AOI221XL U6473 ( .A0(n6416), .A1(n5807), .B0(n6415), .B1(n5806), .C0(n6027), 
        .Y(n5808) );
  INVXL U6474 ( .A(n7317), .Y(n8491) );
  INVXL U6475 ( .A(n8069), .Y(n6891) );
  AOI22XL U6476 ( .A0(n6127), .A1(n6421), .B0(n6126), .B1(n6420), .Y(n7507) );
  AOI21XL U6477 ( .A0(n6415), .A1(n6173), .B0(n6172), .Y(n8340) );
  INVXL U6478 ( .A(n8447), .Y(n8341) );
  INVXL U6479 ( .A(n7570), .Y(n7035) );
  AOI22XL U6480 ( .A0(N2755), .A1(n6418), .B0(N2779), .B1(n6417), .Y(n6419) );
  CLKINVX2 U6481 ( .A(n8070), .Y(n8334) );
  AOI21XL U6482 ( .A0(n3410), .A1(n6872), .B0(n6822), .Y(n6823) );
  AOI21XL U6483 ( .A0(n6821), .A1(n6824), .B0(n3363), .Y(n6822) );
  INVXL U6484 ( .A(n7016), .Y(n6821) );
  INVX4 U6485 ( .A(n3464), .Y(n8496) );
  CLKINVX2 U6486 ( .A(n8419), .Y(n8437) );
  CLKINVX3 U6487 ( .A(n8440), .Y(n8377) );
  CLKINVX2 U6488 ( .A(n7046), .Y(n8441) );
  NOR3X2 U6489 ( .A(n8438), .B(n7046), .C(n7044), .Y(n8444) );
  OAI221XL U6490 ( .A0(op2[0]), .A1(n8466), .B0(n8529), .B1(n8473), .C0(n6313), 
        .Y(n8482) );
  NOR2XL U6491 ( .A(n6401), .B(n6303), .Y(n6317) );
  NOR2XL U6492 ( .A(n6801), .B(n6319), .Y(n6385) );
  AOI211XL U6493 ( .A0(n6303), .A1(n6401), .B0(n6317), .C0(n6299), .Y(n6316)
         );
  INVXL U6494 ( .A(cmd_valid), .Y(n6388) );
  NAND4XL U6495 ( .A(n5486), .B(n5485), .C(n5484), .D(n5483), .Y(n5502) );
  NAND4XL U6496 ( .A(n5402), .B(n5401), .C(n5400), .D(n5399), .Y(n5418) );
  NAND4XL U6497 ( .A(n4540), .B(n4539), .C(n4538), .D(n4537), .Y(n4564) );
  NAND4XL U6498 ( .A(n5528), .B(n5527), .C(n5526), .D(n5525), .Y(n5544) );
  NAND4XL U6499 ( .A(n5444), .B(n5443), .C(n5442), .D(n5441), .Y(n5460) );
  NAND4XL U6500 ( .A(n5360), .B(n5359), .C(n5358), .D(n5357), .Y(n5376) );
  NAND4XL U6501 ( .A(n5318), .B(n5317), .C(n5316), .D(n5315), .Y(n5334) );
  NAND4XL U6502 ( .A(n5276), .B(n5275), .C(n5274), .D(n5273), .Y(n5292) );
  OAI31XL U6503 ( .A0(op2[1]), .A1(n8473), .A2(n8485), .B0(op2[2]), .Y(n8474)
         );
  OAI2BB1XL U6504 ( .A0N(n8527), .A1N(n8486), .B0(n8479), .Y(n3331) );
  AOI211XL U6505 ( .A0(op4[3]), .A1(n6387), .B0(n6386), .C0(n6385), .Y(n3326)
         );
  OAI211XL U6506 ( .A0(n6316), .A1(n8525), .B0(n6306), .C0(n6305), .Y(n3342)
         );
  INVXL U6507 ( .A(n6381), .Y(n3332) );
  AOI22XL U6508 ( .A0(IROM_A[5]), .A1(n8479), .B0(n6382), .B1(n8521), .Y(n3330) );
  AOI21XL U6509 ( .A0(n6323), .A1(n8463), .B0(n6322), .Y(n3328) );
  AOI211XL U6510 ( .A0(n8084), .A1(image_data[0]), .B0(n8083), .C0(n8082), .Y(
        n2808) );
  OAI22XL U6511 ( .A0(n3385), .A1(n8370), .B0(n8323), .B1(n8111), .Y(n8082) );
  AOI21XL U6512 ( .A0(n3367), .A1(n8081), .B0(n8084), .Y(n8083) );
  AOI22XL U6513 ( .A0(n3373), .A1(n8080), .B0(n8417), .B1(n3360), .Y(n8081) );
  AOI211XL U6514 ( .A0(n3351), .A1(n8188), .B0(n7121), .C0(n7120), .Y(n2809)
         );
  AOI2BB2XL U6515 ( .B0(n3346), .B1(n8185), .A0N(n8185), .A1N(image_data[1]), 
        .Y(n7120) );
  AOI22XL U6516 ( .A0(n8438), .A1(n7298), .B0(n8417), .B1(n3375), .Y(n7119) );
  AOI211XL U6517 ( .A0(n7795), .A1(n8188), .B0(n7822), .C0(n7821), .Y(n2810)
         );
  AOI2BB2XL U6518 ( .B0(n3348), .B1(n8185), .A0N(n8185), .A1N(image_data[2]), 
        .Y(n7821) );
  AOI22XL U6519 ( .A0(n8182), .A1(n6880), .B0(n8417), .B1(n3395), .Y(n7820) );
  AOI211XL U6520 ( .A0(n3387), .A1(n8188), .B0(n8187), .C0(n8186), .Y(n2811)
         );
  AOI2BB2XL U6521 ( .B0(n3347), .B1(n8185), .A0N(n8185), .A1N(image_data[3]), 
        .Y(n8186) );
  AOI22XL U6522 ( .A0(n8438), .A1(n3389), .B0(n8182), .B1(n6291), .Y(n8183) );
  AOI211XL U6523 ( .A0(n8503), .A1(n8188), .B0(n7373), .C0(n7372), .Y(n2812)
         );
  AOI2BB2XL U6524 ( .B0(n6855), .B1(n8185), .A0N(n8185), .A1N(image_data[4]), 
        .Y(n7372) );
  AOI22XL U6525 ( .A0(n8417), .A1(n3388), .B0(n8182), .B1(n7326), .Y(n7371) );
  AOI211XL U6526 ( .A0(n3361), .A1(n8188), .B0(n7136), .C0(n7135), .Y(n2813)
         );
  AOI2BB2XL U6527 ( .B0(n7303), .B1(n8185), .A0N(n8185), .A1N(image_data[5]), 
        .Y(n7135) );
  AOI22XL U6528 ( .A0(n8438), .A1(n3357), .B0(n8182), .B1(n7078), .Y(n7134) );
  AOI211XL U6529 ( .A0(n3352), .A1(n8188), .B0(n7658), .C0(n7657), .Y(n2814)
         );
  AOI2BB2XL U6530 ( .B0(n3345), .B1(n8185), .A0N(n8185), .A1N(image_data[6]), 
        .Y(n7657) );
  AOI22XL U6531 ( .A0(n8438), .A1(n3353), .B0(n8417), .B1(n7581), .Y(n7656) );
  AOI211XL U6532 ( .A0(n3362), .A1(n8188), .B0(n6624), .C0(n6623), .Y(n2815)
         );
  AOI2BB2XL U6533 ( .B0(n6959), .B1(n8185), .A0N(n8185), .A1N(image_data[7]), 
        .Y(n6623) );
  AOI22XL U6534 ( .A0(n8438), .A1(n3354), .B0(n8182), .B1(n6651), .Y(n6622) );
  AOI211XL U6535 ( .A0(n3373), .A1(n8099), .B0(n8098), .C0(n8097), .Y(n2816)
         );
  AOI2BB2XL U6536 ( .B0(n3367), .B1(n8096), .A0N(n8096), .A1N(image_data[8]), 
        .Y(n8097) );
  AOI22XL U6537 ( .A0(n8182), .A1(n8114), .B0(n8513), .B1(n3356), .Y(n8095) );
  AOI211XL U6538 ( .A0(n3351), .A1(n8099), .B0(n8006), .C0(n8005), .Y(n2817)
         );
  AOI2BB2XL U6539 ( .B0(n3366), .B1(n8096), .A0N(n8096), .A1N(image_data[9]), 
        .Y(n8005) );
  AOI22XL U6540 ( .A0(n8368), .A1(n3375), .B0(n8513), .B1(n6332), .Y(n8004) );
  AOI211XL U6541 ( .A0(n7795), .A1(n8099), .B0(n7757), .C0(n7756), .Y(n2818)
         );
  AOI2BB2XL U6542 ( .B0(n3348), .B1(n8096), .A0N(n8096), .A1N(image_data[10]), 
        .Y(n7756) );
  AOI22XL U6543 ( .A0(n8513), .A1(n6880), .B0(n8368), .B1(n3395), .Y(n7755) );
  AOI211XL U6544 ( .A0(n3415), .A1(image_data[11]), .B0(n8374), .C0(n8373), 
        .Y(n2819) );
  OAI22XL U6545 ( .A0(n8372), .A1(n8371), .B0(n6407), .B1(n8370), .Y(n8373) );
  AOI21XL U6546 ( .A0(n3347), .A1(n8369), .B0(n3415), .Y(n8374) );
  AOI22XL U6547 ( .A0(n8513), .A1(n6291), .B0(n8368), .B1(n3349), .Y(n8369) );
  AOI211XL U6548 ( .A0(n8503), .A1(n8099), .B0(n8044), .C0(n8043), .Y(n2820)
         );
  AOI2BB2XL U6549 ( .B0(n6855), .B1(n8096), .A0N(n8096), .A1N(image_data[12]), 
        .Y(n8043) );
  AOI22XL U6550 ( .A0(n3371), .A1(n8182), .B0(n8368), .B1(n3388), .Y(n8042) );
  AOI21XL U6551 ( .A0(n3357), .A1(n8182), .B0(n6023), .Y(n2821) );
  OAI221XL U6552 ( .A0(n3415), .A1(n6022), .B0(n8096), .B1(n8552), .C0(n6021), 
        .Y(n6023) );
  AOI22XL U6553 ( .A0(n8368), .A1(n6979), .B0(n8513), .B1(n7078), .Y(n6021) );
  AOI211XL U6554 ( .A0(n3352), .A1(n8099), .B0(n7588), .C0(n7587), .Y(n2822)
         );
  AOI2BB2XL U6555 ( .B0(n3365), .B1(n8096), .A0N(n8096), .A1N(image_data[14]), 
        .Y(n7587) );
  AOI22XL U6556 ( .A0(n8182), .A1(n3353), .B0(n8513), .B1(n3350), .Y(n7586) );
  AOI211XL U6557 ( .A0(n3415), .A1(image_data[15]), .B0(n6972), .C0(n6971), 
        .Y(n2823) );
  OAI22XL U6558 ( .A0(n3394), .A1(n3399), .B0(n7578), .B1(n8371), .Y(n6971) );
  AOI21XL U6559 ( .A0(n6959), .A1(n6969), .B0(n3415), .Y(n6972) );
  AOI22XL U6560 ( .A0(n3354), .A1(n8182), .B0(n8513), .B1(n7035), .Y(n6969) );
  AOI211XL U6561 ( .A0(n3373), .A1(n8416), .B0(n8103), .C0(n8102), .Y(n2824)
         );
  AOI2BB2XL U6562 ( .B0(n3367), .B1(n8413), .A0N(n8413), .A1N(image_data[16]), 
        .Y(n8102) );
  AOI22XL U6563 ( .A0(n8513), .A1(n8114), .B0(n8511), .B1(n3356), .Y(n8100) );
  AOI211XL U6564 ( .A0(n3351), .A1(n8416), .B0(n8003), .C0(n8002), .Y(n2825)
         );
  AOI2BB2XL U6565 ( .B0(n3346), .B1(n8413), .A0N(n8413), .A1N(image_data[17]), 
        .Y(n8002) );
  AOI22XL U6566 ( .A0(n7191), .A1(n8513), .B0(n8512), .B1(n3375), .Y(n8001) );
  AOI211XL U6567 ( .A0(n7795), .A1(n8416), .B0(n7782), .C0(n7781), .Y(n2826)
         );
  AOI2BB2XL U6568 ( .B0(n3348), .B1(n8413), .A0N(n8413), .A1N(image_data[18]), 
        .Y(n7781) );
  AOI22XL U6569 ( .A0(n3358), .A1(n8513), .B0(n8512), .B1(n3395), .Y(n7780) );
  AOI211XL U6570 ( .A0(n3369), .A1(n8416), .B0(n8415), .C0(n8414), .Y(n2827)
         );
  AOI2BB2XL U6571 ( .B0(n3347), .B1(n8413), .A0N(n8413), .A1N(image_data[19]), 
        .Y(n8414) );
  AOI22XL U6572 ( .A0(n3389), .A1(n8513), .B0(n8512), .B1(n3349), .Y(n8411) );
  AOI211XL U6573 ( .A0(n8503), .A1(n8416), .B0(n8061), .C0(n8060), .Y(n2828)
         );
  AOI2BB2XL U6574 ( .B0(n6855), .B1(n8413), .A0N(n8413), .A1N(image_data[20]), 
        .Y(n8060) );
  AOI22XL U6575 ( .A0(n8512), .A1(n3388), .B0(n8511), .B1(n7326), .Y(n8058) );
  AOI211XL U6576 ( .A0(n3361), .A1(n8416), .B0(n7961), .C0(n7960), .Y(n2829)
         );
  AOI2BB2XL U6577 ( .B0(n8496), .B1(n8413), .A0N(n8413), .A1N(image_data[21]), 
        .Y(n7960) );
  AOI22XL U6578 ( .A0(n8512), .A1(n6979), .B0(n8511), .B1(n7078), .Y(n7959) );
  AOI22XL U6579 ( .A0(n8513), .A1(n3353), .B0(n8512), .B1(n7581), .Y(n8514) );
  AOI21XL U6580 ( .A0(n8511), .A1(n3350), .B0(n8510), .Y(n8515) );
  AOI211XL U6581 ( .A0(n3362), .A1(n8416), .B0(n7038), .C0(n7037), .Y(n2831)
         );
  AOI2BB2XL U6582 ( .B0(n6959), .B1(n8413), .A0N(n8413), .A1N(image_data[23]), 
        .Y(n7037) );
  AOI22XL U6583 ( .A0(n3354), .A1(n8513), .B0(n8511), .B1(n7035), .Y(n7036) );
  AOI211XL U6584 ( .A0(n3355), .A1(n8451), .B0(n8123), .C0(n8122), .Y(n2832)
         );
  AOI2BB2XL U6585 ( .B0(n3367), .B1(n8448), .A0N(n8448), .A1N(image_data[24]), 
        .Y(n8122) );
  AOI22XL U6586 ( .A0(n6145), .A1(n8511), .B0(n3379), .B1(n3360), .Y(n8121) );
  AOI211XL U6587 ( .A0(n3351), .A1(n8451), .B0(n8016), .C0(n8015), .Y(n2833)
         );
  AOI2BB2XL U6588 ( .B0(n3366), .B1(n8448), .A0N(n8448), .A1N(image_data[25]), 
        .Y(n8015) );
  AOI22XL U6589 ( .A0(n7298), .A1(n8511), .B0(n3379), .B1(n3375), .Y(n8013) );
  AOI211XL U6590 ( .A0(n7795), .A1(n8451), .B0(n7785), .C0(n7784), .Y(n2834)
         );
  AOI2BB2XL U6591 ( .B0(n3348), .B1(n8448), .A0N(n8448), .A1N(image_data[26]), 
        .Y(n7784) );
  AOI22XL U6592 ( .A0(n8032), .A1(n6880), .B0(n3379), .B1(n3395), .Y(n7783) );
  AOI211XL U6593 ( .A0(n3369), .A1(n8451), .B0(n8450), .C0(n8449), .Y(n2835)
         );
  AOI2BB2XL U6594 ( .B0(n3347), .B1(n8448), .A0N(n8448), .A1N(image_data[27]), 
        .Y(n8449) );
  AOI22XL U6595 ( .A0(n3389), .A1(n8511), .B0(n3379), .B1(n3349), .Y(n8445) );
  AOI211XL U6596 ( .A0(n8451), .A1(n8503), .B0(n8037), .C0(n8036), .Y(n2836)
         );
  OAI2BB2XL U6597 ( .B0(n8035), .B1(n8412), .A0N(n8034), .A1N(image_data[28]), 
        .Y(n8036) );
  AOI21XL U6598 ( .A0(n6855), .A1(n8033), .B0(n8034), .Y(n8037) );
  AOI22XL U6599 ( .A0(n3379), .A1(n3388), .B0(n8032), .B1(n7326), .Y(n8033) );
  AOI211XL U6600 ( .A0(n3361), .A1(n8451), .B0(n7971), .C0(n7970), .Y(n2837)
         );
  AOI2BB2XL U6601 ( .B0(n8496), .B1(n8448), .A0N(n8448), .A1N(image_data[29]), 
        .Y(n7970) );
  AOI22XL U6602 ( .A0(n3379), .A1(n6979), .B0(n8032), .B1(n7078), .Y(n7969) );
  AOI21XL U6603 ( .A0(n3352), .A1(n8451), .B0(n5906), .Y(n2838) );
  AOI22XL U6604 ( .A0(n8511), .A1(n3353), .B0(n3379), .B1(n7581), .Y(n5904) );
  AOI211XL U6605 ( .A0(n3362), .A1(n8451), .B0(n7051), .C0(n7050), .Y(n2839)
         );
  AOI2BB2XL U6606 ( .B0(n6959), .B1(n8448), .A0N(n8448), .A1N(image_data[31]), 
        .Y(n7050) );
  AOI22XL U6607 ( .A0(n8032), .A1(n6651), .B0(n3379), .B1(n3368), .Y(n7049) );
  AOI211XL U6608 ( .A0(n3355), .A1(n8403), .B0(n8109), .C0(n8108), .Y(n2840)
         );
  AOI2BB2XL U6609 ( .B0(n3367), .B1(n8400), .A0N(n8400), .A1N(image_data[32]), 
        .Y(n8108) );
  AOI22XL U6610 ( .A0(n3376), .A1(n3356), .B0(n8398), .B1(n3360), .Y(n8107) );
  AOI211XL U6611 ( .A0(n3351), .A1(n8403), .B0(n7990), .C0(n7989), .Y(n2841)
         );
  AOI2BB2XL U6612 ( .B0(n3366), .B1(n8400), .A0N(n8400), .A1N(image_data[33]), 
        .Y(n7989) );
  AOI22XL U6613 ( .A0(n3376), .A1(n6332), .B0(n8398), .B1(n3375), .Y(n7988) );
  AOI211XL U6614 ( .A0(n7795), .A1(n8403), .B0(n7764), .C0(n7763), .Y(n2842)
         );
  AOI2BB2XL U6615 ( .B0(n3348), .B1(n8400), .A0N(n8400), .A1N(image_data[34]), 
        .Y(n7763) );
  AOI22XL U6616 ( .A0(n3376), .A1(n6880), .B0(n8398), .B1(n7761), .Y(n7762) );
  AOI211XL U6617 ( .A0(n3369), .A1(n8403), .B0(n8402), .C0(n8401), .Y(n2843)
         );
  AOI2BB2XL U6618 ( .B0(n3347), .B1(n8400), .A0N(n8400), .A1N(image_data[35]), 
        .Y(n8401) );
  AOI22XL U6619 ( .A0(n3376), .A1(n6291), .B0(n8398), .B1(n3349), .Y(n8399) );
  AOI211XL U6620 ( .A0(n8503), .A1(n8403), .B0(n8050), .C0(n8049), .Y(n2844)
         );
  AOI2BB2XL U6621 ( .B0(n6855), .B1(n8400), .A0N(n8400), .A1N(image_data[36]), 
        .Y(n8049) );
  AOI22XL U6622 ( .A0(n3376), .A1(n7326), .B0(n8398), .B1(n3388), .Y(n8048) );
  AOI211XL U6623 ( .A0(n3361), .A1(n8403), .B0(n7948), .C0(n7947), .Y(n2845)
         );
  AOI2BB2XL U6624 ( .B0(n8496), .B1(n8400), .A0N(n8400), .A1N(image_data[37]), 
        .Y(n7947) );
  AOI22XL U6625 ( .A0(n3376), .A1(n7078), .B0(n8398), .B1(n6979), .Y(n7946) );
  AOI211XL U6626 ( .A0(n3352), .A1(n8403), .B0(n7597), .C0(n7596), .Y(n2846)
         );
  AOI2BB2XL U6627 ( .B0(n3365), .B1(n8400), .A0N(n8400), .A1N(image_data[38]), 
        .Y(n7596) );
  AOI22XL U6628 ( .A0(n3376), .A1(n3350), .B0(n8398), .B1(n7581), .Y(n7595) );
  AOI211XL U6629 ( .A0(n3362), .A1(n8403), .B0(n7013), .C0(n7012), .Y(n2847)
         );
  AOI2BB2XL U6630 ( .B0(n6959), .B1(n8400), .A0N(n8400), .A1N(image_data[39]), 
        .Y(n7012) );
  AOI22XL U6631 ( .A0(n3376), .A1(n6651), .B0(n8398), .B1(n3368), .Y(n7011) );
  AOI211XL U6632 ( .A0(n3355), .A1(n8089), .B0(n8088), .C0(n8087), .Y(n2848)
         );
  AOI2BB2XL U6633 ( .B0(n3367), .B1(n8086), .A0N(n8086), .A1N(image_data[40]), 
        .Y(n8087) );
  AOI22XL U6634 ( .A0(n3376), .A1(n8114), .B0(n8385), .B1(n3360), .Y(n8085) );
  AOI211XL U6635 ( .A0(n3351), .A1(n8089), .B0(n7997), .C0(n7996), .Y(n2849)
         );
  AOI2BB2XL U6636 ( .B0(n3366), .B1(n8086), .A0N(n8086), .A1N(image_data[41]), 
        .Y(n7996) );
  AOI22XL U6637 ( .A0(n8038), .A1(n6332), .B0(n3376), .B1(n7298), .Y(n7994) );
  AOI211XL U6638 ( .A0(n7795), .A1(n8089), .B0(n7753), .C0(n7752), .Y(n2850)
         );
  AOI2BB2XL U6639 ( .B0(n3348), .B1(n8086), .A0N(n8086), .A1N(image_data[42]), 
        .Y(n7752) );
  AOI22XL U6640 ( .A0(n8038), .A1(n6880), .B0(n3376), .B1(n3358), .Y(n7751) );
  AOI21XL U6641 ( .A0(n3376), .A1(n8423), .B0(n6364), .Y(n2851) );
  AOI22XL U6642 ( .A0(n8038), .A1(n6291), .B0(n8385), .B1(n3349), .Y(n6362) );
  AOI211XL U6643 ( .A0(n8503), .A1(n8089), .B0(n8047), .C0(n8046), .Y(n2852)
         );
  AOI2BB2XL U6644 ( .B0(n6855), .B1(n8086), .A0N(n8086), .A1N(image_data[44]), 
        .Y(n8046) );
  AOI22XL U6645 ( .A0(n3376), .A1(n3371), .B0(n8385), .B1(n3388), .Y(n8045) );
  AOI211XL U6646 ( .A0(n3361), .A1(n8089), .B0(n7951), .C0(n7950), .Y(n2853)
         );
  AOI2BB2XL U6647 ( .B0(n8496), .B1(n8086), .A0N(n8086), .A1N(image_data[45]), 
        .Y(n7950) );
  AOI22XL U6648 ( .A0(n3376), .A1(n3357), .B0(n8385), .B1(n6979), .Y(n7949) );
  AOI21XL U6649 ( .A0(n3376), .A1(n3353), .B0(n6358), .Y(n2854) );
  AOI2BB2XL U6650 ( .B0(n6357), .B1(n8086), .A0N(n8086), .A1N(image_data[46]), 
        .Y(n6358) );
  AOI211XL U6651 ( .A0(n6975), .A1(n3352), .B0(n3440), .C0(n6354), .Y(n6357)
         );
  OAI22XL U6652 ( .A0(n3396), .A1(n8432), .B0(n7740), .B1(n7995), .Y(n6354) );
  AOI211XL U6653 ( .A0(n6978), .A1(image_data[47]), .B0(n6977), .C0(n6976), 
        .Y(n2855) );
  OAI22XL U6654 ( .A0(n3394), .A1(n7995), .B0(n7578), .B1(n7750), .Y(n6976) );
  AOI21XL U6655 ( .A0(n6959), .A1(n6974), .B0(n6978), .Y(n6977) );
  AOI22XL U6656 ( .A0(n8038), .A1(n6651), .B0(n3376), .B1(n6973), .Y(n6974) );
  AOI2BB2XL U6657 ( .B0(n3367), .B1(n8433), .A0N(n8433), .A1N(image_data[48]), 
        .Y(n8112) );
  AOI22XL U6658 ( .A0(n8430), .A1(n3360), .B0(n8437), .B1(n3356), .Y(n8110) );
  AOI211XL U6659 ( .A0(n3351), .A1(n8436), .B0(n8009), .C0(n8008), .Y(n2857)
         );
  AOI2BB2XL U6660 ( .B0(n3346), .B1(n8433), .A0N(n8433), .A1N(image_data[49]), 
        .Y(n8008) );
  AOI22XL U6661 ( .A0(n8430), .A1(n3375), .B0(n8437), .B1(n6332), .Y(n8007) );
  AOI211XL U6662 ( .A0(n8436), .A1(n7795), .B0(n7749), .C0(n7748), .Y(n2858)
         );
  OAI2BB2XL U6663 ( .B0(n3372), .B1(n8454), .A0N(image_data[50]), .A1N(n7747), 
        .Y(n7748) );
  AOI21XL U6664 ( .A0(n3348), .A1(n7746), .B0(n7747), .Y(n7749) );
  AOI22XL U6665 ( .A0(n8038), .A1(n3358), .B0(n8437), .B1(n6880), .Y(n7746) );
  AOI2BB2XL U6666 ( .B0(n3347), .B1(n8433), .A0N(n8433), .A1N(image_data[51]), 
        .Y(n8434) );
  AOI22XL U6667 ( .A0(n8437), .A1(n6291), .B0(n8430), .B1(n3349), .Y(n8431) );
  AOI211XL U6668 ( .A0(n8503), .A1(n8436), .B0(n8041), .C0(n8040), .Y(n2860)
         );
  AOI2BB2XL U6669 ( .B0(n6855), .B1(n8433), .A0N(n8433), .A1N(image_data[52]), 
        .Y(n8040) );
  AOI22XL U6670 ( .A0(n8038), .A1(n3371), .B0(n8430), .B1(n3388), .Y(n8039) );
  AOI211XL U6671 ( .A0(n3361), .A1(n8436), .B0(n7945), .C0(n7944), .Y(n2861)
         );
  AOI2BB2XL U6672 ( .B0(n8496), .B1(n8433), .A0N(n8433), .A1N(image_data[53]), 
        .Y(n7944) );
  AOI22XL U6673 ( .A0(n8038), .A1(n3357), .B0(n8430), .B1(n6979), .Y(n7943) );
  AOI211XL U6674 ( .A0(n3352), .A1(n8436), .B0(n7603), .C0(n7602), .Y(n2862)
         );
  AOI2BB2XL U6675 ( .B0(n3365), .B1(n8433), .A0N(n8433), .A1N(image_data[54]), 
        .Y(n7602) );
  AOI22XL U6676 ( .A0(n8430), .A1(n7581), .B0(n8437), .B1(n3350), .Y(n7601) );
  AOI211XL U6677 ( .A0(n3362), .A1(n8436), .B0(n7019), .C0(n7018), .Y(n2863)
         );
  AOI2BB2XL U6678 ( .B0(n6959), .B1(n8433), .A0N(n8433), .A1N(image_data[55]), 
        .Y(n7018) );
  AOI22XL U6679 ( .A0(n8437), .A1(n6651), .B0(n8430), .B1(n3368), .Y(n7017) );
  AOI211XL U6680 ( .A0(n3373), .A1(n3429), .B0(n8106), .C0(n8105), .Y(n2864)
         );
  AOI2BB2XL U6681 ( .B0(n3367), .B1(n8420), .A0N(n8420), .A1N(image_data[56]), 
        .Y(n8105) );
  AOI22XL U6682 ( .A0(n8452), .A1(n3360), .B0(n8417), .B1(n3356), .Y(n8104) );
  AOI211XL U6683 ( .A0(n3351), .A1(n3429), .B0(n7993), .C0(n7992), .Y(n2865)
         );
  AOI2BB2XL U6684 ( .B0(n3346), .B1(n8420), .A0N(n8420), .A1N(image_data[57]), 
        .Y(n7992) );
  AOI22XL U6685 ( .A0(n8452), .A1(n3375), .B0(n8417), .B1(n6332), .Y(n7991) );
  AOI211XL U6686 ( .A0(n7795), .A1(n3429), .B0(n7776), .C0(n7775), .Y(n2866)
         );
  AOI2BB2XL U6687 ( .B0(n3348), .B1(n8420), .A0N(n8420), .A1N(image_data[58]), 
        .Y(n7775) );
  AOI22XL U6688 ( .A0(n8417), .A1(n6880), .B0(n8452), .B1(n3395), .Y(n7774) );
  AOI211XL U6689 ( .A0(n3369), .A1(n3429), .B0(n8422), .C0(n8421), .Y(n2867)
         );
  AOI2BB2XL U6690 ( .B0(n3347), .B1(n8420), .A0N(n8420), .A1N(image_data[59]), 
        .Y(n8421) );
  AOI22XL U6691 ( .A0(n8417), .A1(n6291), .B0(n8452), .B1(n3349), .Y(n8418) );
  AOI211XL U6692 ( .A0(n8503), .A1(n3429), .B0(n8053), .C0(n8052), .Y(n2868)
         );
  AOI2BB2XL U6693 ( .B0(n6855), .B1(n8420), .A0N(n8420), .A1N(image_data[60]), 
        .Y(n8052) );
  AOI22XL U6694 ( .A0(n8452), .A1(n3388), .B0(n8417), .B1(n7326), .Y(n8051) );
  AOI211XL U6695 ( .A0(n3361), .A1(n3429), .B0(n7954), .C0(n7953), .Y(n2869)
         );
  AOI2BB2XL U6696 ( .B0(n8496), .B1(n8420), .A0N(n8420), .A1N(image_data[61]), 
        .Y(n7953) );
  AOI22XL U6697 ( .A0(n8452), .A1(n6979), .B0(n8417), .B1(n7078), .Y(n7952) );
  AOI211XL U6698 ( .A0(n3352), .A1(n3429), .B0(n7609), .C0(n7608), .Y(n2870)
         );
  AOI2BB2XL U6699 ( .B0(n3365), .B1(n8420), .A0N(n8420), .A1N(image_data[62]), 
        .Y(n7608) );
  AOI22XL U6700 ( .A0(n8452), .A1(n7581), .B0(n8417), .B1(n3350), .Y(n7607) );
  AOI211XL U6701 ( .A0(n3362), .A1(n3429), .B0(n7025), .C0(n7024), .Y(n2871)
         );
  AOI2BB2XL U6702 ( .B0(n6959), .B1(n8420), .A0N(n8420), .A1N(image_data[63]), 
        .Y(n7024) );
  AOI22XL U6703 ( .A0(n8417), .A1(n6651), .B0(n8452), .B1(n3368), .Y(n7022) );
  AOI211XL U6704 ( .A0(n3355), .A1(n8094), .B0(n8093), .C0(n8092), .Y(n2872)
         );
  AOI2BB2XL U6705 ( .B0(n3367), .B1(n8091), .A0N(n8091), .A1N(image_data[64]), 
        .Y(n8092) );
  AOI22XL U6706 ( .A0(n8114), .A1(n8417), .B0(n8200), .B1(n3360), .Y(n8090) );
  AOI211XL U6707 ( .A0(n3351), .A1(n8094), .B0(n8000), .C0(n7999), .Y(n2873)
         );
  AOI2BB2XL U6708 ( .B0(n3366), .B1(n8091), .A0N(n8091), .A1N(image_data[65]), 
        .Y(n7999) );
  AOI22XL U6709 ( .A0(n7298), .A1(n8417), .B0(n8200), .B1(n3375), .Y(n7998) );
  AOI211XL U6710 ( .A0(n7795), .A1(n8094), .B0(n7779), .C0(n7778), .Y(n2874)
         );
  AOI2BB2XL U6711 ( .B0(n3348), .B1(n8091), .A0N(n8091), .A1N(image_data[66]), 
        .Y(n7778) );
  AOI22XL U6712 ( .A0(n3358), .A1(n8417), .B0(n8368), .B1(n6880), .Y(n7777) );
  AOI21XL U6713 ( .A0(n3369), .A1(n8094), .B0(n6270), .Y(n2875) );
  AOI22XL U6714 ( .A0(n8368), .A1(n6291), .B0(n8200), .B1(n3349), .Y(n6267) );
  AOI211XL U6715 ( .A0(n8503), .A1(n8094), .B0(n8057), .C0(n8056), .Y(n2876)
         );
  AOI2BB2XL U6716 ( .B0(n6855), .B1(n8091), .A0N(n8091), .A1N(image_data[68]), 
        .Y(n8056) );
  AOI22XL U6717 ( .A0(n3371), .A1(n8417), .B0(n8200), .B1(n3388), .Y(n8054) );
  AOI211XL U6718 ( .A0(n3361), .A1(n8094), .B0(n7958), .C0(n7957), .Y(n2877)
         );
  AOI2BB2XL U6719 ( .B0(n8496), .B1(n8091), .A0N(n8091), .A1N(image_data[69]), 
        .Y(n7957) );
  AOI22XL U6720 ( .A0(n3357), .A1(n8417), .B0(n8200), .B1(n6979), .Y(n7955) );
  AOI211XL U6721 ( .A0(n3352), .A1(n8094), .B0(n7612), .C0(n7611), .Y(n2878)
         );
  AOI2BB2XL U6722 ( .B0(n3365), .B1(n8091), .A0N(n8091), .A1N(image_data[70]), 
        .Y(n7611) );
  AOI22XL U6723 ( .A0(n8417), .A1(n3353), .B0(n8200), .B1(n7581), .Y(n7610) );
  AOI211XL U6724 ( .A0(n3362), .A1(n8094), .B0(n7028), .C0(n7027), .Y(n2879)
         );
  AOI2BB2XL U6725 ( .B0(n6959), .B1(n8091), .A0N(n8091), .A1N(image_data[71]), 
        .Y(n7027) );
  AOI22XL U6726 ( .A0(n3354), .A1(n8417), .B0(n8368), .B1(n6651), .Y(n7026) );
  AOI22XL U6727 ( .A0(n8260), .A1(n3360), .B0(n8512), .B1(n3356), .Y(n6999) );
  AOI211XL U6728 ( .A0(n3351), .A1(n8031), .B0(n8020), .C0(n8019), .Y(n2881)
         );
  AOI2BB2XL U6729 ( .B0(n3346), .B1(n8018), .A0N(n8018), .A1N(image_data[73]), 
        .Y(n8019) );
  AOI22XL U6730 ( .A0(n8260), .A1(n3375), .B0(n8512), .B1(n6332), .Y(n8017) );
  AOI211XL U6731 ( .A0(n8031), .A1(n7795), .B0(n6949), .C0(n6948), .Y(n2882)
         );
  NOR2XL U6732 ( .A(n7773), .B(n3399), .Y(n6949) );
  AOI22XL U6733 ( .A0(n8512), .A1(n6880), .B0(n8260), .B1(n3395), .Y(n6947) );
  AOI21XL U6734 ( .A0(n3389), .A1(n8368), .B0(n6368), .Y(n2883) );
  AOI2BB2XL U6735 ( .B0(n6367), .B1(n8018), .A0N(n8018), .A1N(image_data[75]), 
        .Y(n6368) );
  AOI211XL U6736 ( .A0(n7582), .A1(n3369), .B0(n6403), .C0(n6365), .Y(n6367)
         );
  OAI22XL U6737 ( .A0(n8447), .A1(n8101), .B0(n3386), .B1(n7684), .Y(n6365) );
  AOI211XL U6738 ( .A0(n8031), .A1(n8503), .B0(n8030), .C0(n8029), .Y(n2884)
         );
  OAI2BB2XL U6739 ( .B0(n8055), .B1(n8101), .A0N(image_data[76]), .A1N(n3454), 
        .Y(n8029) );
  AOI22XL U6740 ( .A0(n3371), .A1(n8368), .B0(n8260), .B1(n3388), .Y(n8027) );
  AOI211XL U6741 ( .A0(n8031), .A1(n3361), .B0(n7057), .C0(n7056), .Y(n2885)
         );
  NOR2XL U6742 ( .A(n3391), .B(n3399), .Y(n7057) );
  AOI22XL U6743 ( .A0(n8260), .A1(n6979), .B0(n8512), .B1(n7078), .Y(n7055) );
  OAI22XL U6744 ( .A0(n3396), .A1(n8101), .B0(n3399), .B1(n3392), .Y(n7584) );
  AOI22XL U6745 ( .A0(n3352), .A1(n7582), .B0(n8260), .B1(n7581), .Y(n7583) );
  AOI211XL U6746 ( .A0(n3362), .A1(n8031), .B0(n7054), .C0(n7053), .Y(n2887)
         );
  AOI2BB2XL U6747 ( .B0(n6959), .B1(n8018), .A0N(n8018), .A1N(image_data[79]), 
        .Y(n7053) );
  AOI22XL U6748 ( .A0(n3354), .A1(n8368), .B0(n8512), .B1(n6651), .Y(n7052) );
  AOI211XL U6749 ( .A0(n3355), .A1(n8429), .B0(n8117), .C0(n8116), .Y(n2888)
         );
  AOI2BB2XL U6750 ( .B0(n3367), .B1(n8426), .A0N(n8426), .A1N(image_data[80]), 
        .Y(n8116) );
  AOI22XL U6751 ( .A0(n8512), .A1(n8114), .B0(n3379), .B1(n3356), .Y(n8115) );
  AOI211XL U6752 ( .A0(n3351), .A1(n8429), .B0(n7233), .C0(n7232), .Y(n2889)
         );
  AOI2BB2XL U6753 ( .B0(n3346), .B1(n8426), .A0N(n8426), .A1N(image_data[81]), 
        .Y(n7232) );
  AOI22XL U6754 ( .A0(n8512), .A1(n7298), .B0(n3379), .B1(n6332), .Y(n7231) );
  AOI21XL U6755 ( .A0(n6879), .A1(n8429), .B0(n5272), .Y(n2890) );
  AOI22XL U6756 ( .A0(n3358), .A1(n8512), .B0(n3379), .B1(n6880), .Y(n5270) );
  AOI211XL U6757 ( .A0(n3369), .A1(n8429), .B0(n8428), .C0(n8427), .Y(n2891)
         );
  AOI2BB2XL U6758 ( .B0(n3347), .B1(n8426), .A0N(n8426), .A1N(image_data[83]), 
        .Y(n8427) );
  AOI22XL U6759 ( .A0(n8423), .A1(n8512), .B0(n3379), .B1(n6291), .Y(n8424) );
  AOI211XL U6760 ( .A0(n8503), .A1(n8429), .B0(n8064), .C0(n8063), .Y(n2892)
         );
  AOI2BB2XL U6761 ( .B0(n6855), .B1(n8426), .A0N(n8426), .A1N(image_data[84]), 
        .Y(n8063) );
  AOI22XL U6762 ( .A0(n3371), .A1(n8512), .B0(n3379), .B1(n7326), .Y(n8062) );
  AOI211XL U6763 ( .A0(n3361), .A1(n8429), .B0(n7965), .C0(n7964), .Y(n2893)
         );
  AOI2BB2XL U6764 ( .B0(n8496), .B1(n8426), .A0N(n8426), .A1N(image_data[85]), 
        .Y(n7964) );
  AOI22XL U6765 ( .A0(n3357), .A1(n8512), .B0(n3379), .B1(n7078), .Y(n7962) );
  AOI211XL U6766 ( .A0(n3352), .A1(n8429), .B0(n7615), .C0(n7614), .Y(n2894)
         );
  AOI2BB2XL U6767 ( .B0(n3365), .B1(n8426), .A0N(n8426), .A1N(image_data[86]), 
        .Y(n7614) );
  AOI22XL U6768 ( .A0(n8512), .A1(n3353), .B0(n3379), .B1(n3350), .Y(n7613) );
  AOI221XL U6769 ( .A0(image_data[87]), .A1(n7564), .B0(n7563), .B1(n8426), 
        .C0(n7562), .Y(n2895) );
  AOI22XL U6770 ( .A0(n3379), .A1(n6651), .B0(n8259), .B1(n3368), .Y(n7561) );
  AOI211XL U6771 ( .A0(n3373), .A1(n8410), .B0(n7370), .C0(n7369), .Y(n2896)
         );
  AOI2BB2XL U6772 ( .B0(n3344), .B1(n8407), .A0N(n8407), .A1N(image_data[88]), 
        .Y(n7369) );
  AOI22XL U6773 ( .A0(n8114), .A1(n3379), .B0(n8404), .B1(n3360), .Y(n7368) );
  AOI211XL U6774 ( .A0(n3351), .A1(n8410), .B0(n7100), .C0(n7099), .Y(n2897)
         );
  AOI2BB2XL U6775 ( .B0(n3366), .B1(n8407), .A0N(n8407), .A1N(image_data[89]), 
        .Y(n7099) );
  AOI22XL U6776 ( .A0(n7298), .A1(n3379), .B0(n8404), .B1(n3375), .Y(n7098) );
  AOI211XL U6777 ( .A0(n7795), .A1(n8410), .B0(n7760), .C0(n7759), .Y(n2898)
         );
  AOI2BB2XL U6778 ( .B0(n3348), .B1(n8407), .A0N(n8407), .A1N(image_data[90]), 
        .Y(n7759) );
  AOI22XL U6779 ( .A0(n3358), .A1(n3379), .B0(n8404), .B1(n3395), .Y(n7758) );
  AOI211XL U6780 ( .A0(n3369), .A1(n8410), .B0(n8409), .C0(n8408), .Y(n2899)
         );
  AOI2BB2XL U6781 ( .B0(n3347), .B1(n8407), .A0N(n8407), .A1N(image_data[91]), 
        .Y(n8408) );
  AOI22XL U6782 ( .A0(n8423), .A1(n3379), .B0(n8404), .B1(n3349), .Y(n8405) );
  AOI211XL U6783 ( .A0(n8503), .A1(n8410), .B0(n7367), .C0(n7366), .Y(n2900)
         );
  AOI2BB2XL U6784 ( .B0(n6855), .B1(n8407), .A0N(n8407), .A1N(image_data[92]), 
        .Y(n7366) );
  AOI22XL U6785 ( .A0(n3371), .A1(n3379), .B0(n8404), .B1(n3388), .Y(n7365) );
  AOI211XL U6786 ( .A0(n3361), .A1(n8410), .B0(n7103), .C0(n7102), .Y(n2901)
         );
  AOI2BB2XL U6787 ( .B0(n8496), .B1(n8407), .A0N(n8407), .A1N(image_data[93]), 
        .Y(n7102) );
  AOI22XL U6788 ( .A0(n3357), .A1(n3379), .B0(n8404), .B1(n6979), .Y(n7101) );
  AOI211XL U6789 ( .A0(n3352), .A1(n8410), .B0(n7591), .C0(n7590), .Y(n2902)
         );
  AOI2BB2XL U6790 ( .B0(n3365), .B1(n8407), .A0N(n8407), .A1N(image_data[94]), 
        .Y(n7590) );
  AOI22XL U6791 ( .A0(n3379), .A1(n3353), .B0(n8404), .B1(n7581), .Y(n7589) );
  AOI221XL U6792 ( .A0(image_data[95]), .A1(n7575), .B0(n7574), .B1(n8407), 
        .C0(n7573), .Y(n2903) );
  AOI22XL U6793 ( .A0(n3354), .A1(n3379), .B0(n8404), .B1(n3368), .Y(n7571) );
  AOI211XL U6794 ( .A0(n3355), .A1(n7769), .B0(n7437), .C0(n7436), .Y(n2904)
         );
  AOI2BB2XL U6795 ( .B0(n3344), .B1(n7766), .A0N(n7766), .A1N(image_data[96]), 
        .Y(n7436) );
  AOI22XL U6796 ( .A0(n8114), .A1(n8398), .B0(n8207), .B1(n3360), .Y(n7435) );
  AOI211XL U6797 ( .A0(n3351), .A1(n7769), .B0(n7190), .C0(n7189), .Y(n2905)
         );
  AOI2BB2XL U6798 ( .B0(n3346), .B1(n7766), .A0N(n7766), .A1N(image_data[97]), 
        .Y(n7189) );
  AOI22XL U6799 ( .A0(n7191), .A1(n8398), .B0(n8207), .B1(n3375), .Y(n7188) );
  AOI211XL U6800 ( .A0(n7795), .A1(n7769), .B0(n7768), .C0(n7767), .Y(n2906)
         );
  AOI2BB2XL U6801 ( .B0(n3348), .B1(n7766), .A0N(n7766), .A1N(image_data[98]), 
        .Y(n7767) );
  AOI22XL U6802 ( .A0(n3358), .A1(n8398), .B0(n8207), .B1(n3395), .Y(n7765) );
  AOI221XL U6803 ( .A0(image_data[99]), .A1(n7003), .B0(n6410), .B1(n7766), 
        .C0(n6409), .Y(n2907) );
  AOI22XL U6804 ( .A0(n8385), .A1(n6291), .B0(n8207), .B1(n3349), .Y(n6408) );
  AOI211XL U6805 ( .A0(n8503), .A1(n7769), .B0(n7440), .C0(n7439), .Y(n2908)
         );
  AOI2BB2XL U6806 ( .B0(n6855), .B1(n7766), .A0N(n7766), .A1N(image_data[100]), 
        .Y(n7439) );
  AOI22XL U6807 ( .A0(n3371), .A1(n8398), .B0(n8207), .B1(n3388), .Y(n7438) );
  AOI211XL U6808 ( .A0(n3361), .A1(n7769), .B0(n7187), .C0(n7186), .Y(n2909)
         );
  AOI2BB2XL U6809 ( .B0(n8496), .B1(n7766), .A0N(n7766), .A1N(image_data[101]), 
        .Y(n7186) );
  AOI22XL U6810 ( .A0(n3357), .A1(n8398), .B0(n8207), .B1(n6979), .Y(n7185) );
  AOI211XL U6811 ( .A0(n3352), .A1(n7769), .B0(n7600), .C0(n7599), .Y(n2910)
         );
  AOI2BB2XL U6812 ( .B0(n3365), .B1(n7766), .A0N(n7766), .A1N(image_data[102]), 
        .Y(n7599) );
  AOI22XL U6813 ( .A0(n8398), .A1(n3353), .B0(n8207), .B1(n7581), .Y(n7598) );
  AOI211XL U6814 ( .A0(n3362), .A1(n7769), .B0(n7006), .C0(n7005), .Y(n2911)
         );
  AOI2BB2XL U6815 ( .B0(n6959), .B1(n7766), .A0N(n7766), .A1N(image_data[103]), 
        .Y(n7005) );
  AOI22XL U6816 ( .A0(n3354), .A1(n8398), .B0(n8207), .B1(n3368), .Y(n7004) );
  AOI211XL U6817 ( .A0(n3355), .A1(n8391), .B0(n7460), .C0(n7459), .Y(n2912)
         );
  AOI2BB2XL U6818 ( .B0(n3344), .B1(n8388), .A0N(n8388), .A1N(image_data[104]), 
        .Y(n7459) );
  AOI22XL U6819 ( .A0(n8385), .A1(n8114), .B0(n8430), .B1(n3356), .Y(n7458) );
  AOI211XL U6820 ( .A0(n3351), .A1(n8391), .B0(n7212), .C0(n7211), .Y(n2913)
         );
  AOI2BB2XL U6821 ( .B0(n3346), .B1(n8388), .A0N(n8388), .A1N(image_data[105]), 
        .Y(n7211) );
  AOI22XL U6822 ( .A0(n8385), .A1(n7298), .B0(n8430), .B1(n6332), .Y(n7210) );
  AOI211XL U6823 ( .A0(n7795), .A1(n8391), .B0(n7772), .C0(n7771), .Y(n2914)
         );
  AOI2BB2XL U6824 ( .B0(n3348), .B1(n8388), .A0N(n8388), .A1N(image_data[106]), 
        .Y(n7771) );
  AOI22XL U6825 ( .A0(n3358), .A1(n8385), .B0(n8430), .B1(n6880), .Y(n7770) );
  AOI211XL U6826 ( .A0(n3369), .A1(n8391), .B0(n8390), .C0(n8389), .Y(n2915)
         );
  AOI2BB2XL U6827 ( .B0(n3347), .B1(n8388), .A0N(n8388), .A1N(image_data[107]), 
        .Y(n8389) );
  AOI22XL U6828 ( .A0(n8423), .A1(n8385), .B0(n8430), .B1(n6291), .Y(n8386) );
  AOI211XL U6829 ( .A0(n8503), .A1(n8391), .B0(n7466), .C0(n7465), .Y(n2916)
         );
  AOI2BB2XL U6830 ( .B0(n6855), .B1(n8388), .A0N(n8388), .A1N(image_data[108]), 
        .Y(n7465) );
  AOI22XL U6831 ( .A0(n3371), .A1(n8385), .B0(n8430), .B1(n7326), .Y(n7464) );
  AOI211XL U6832 ( .A0(n3361), .A1(n8391), .B0(n7221), .C0(n7220), .Y(n2917)
         );
  AOI2BB2XL U6833 ( .B0(n8496), .B1(n8388), .A0N(n8388), .A1N(image_data[109]), 
        .Y(n7220) );
  AOI22XL U6834 ( .A0(n3357), .A1(n8385), .B0(n8430), .B1(n7078), .Y(n7219) );
  AOI211XL U6835 ( .A0(n3352), .A1(n8391), .B0(n7606), .C0(n7605), .Y(n2918)
         );
  AOI2BB2XL U6836 ( .B0(n3365), .B1(n8388), .A0N(n8388), .A1N(image_data[110]), 
        .Y(n7605) );
  AOI22XL U6837 ( .A0(n8385), .A1(n3353), .B0(n8430), .B1(n3350), .Y(n7604) );
  AOI211XL U6838 ( .A0(n3362), .A1(n8391), .B0(n6709), .C0(n6708), .Y(n2919)
         );
  AOI2BB2XL U6839 ( .B0(n6586), .B1(n8388), .A0N(n8388), .A1N(image_data[111]), 
        .Y(n6708) );
  AOI22XL U6840 ( .A0(n3354), .A1(n8385), .B0(n8430), .B1(n6651), .Y(n6706) );
  AOI211XL U6841 ( .A0(n3355), .A1(n3428), .B0(n7541), .C0(n7540), .Y(n2920)
         );
  AOI2BB2XL U6842 ( .B0(n3367), .B1(n8455), .A0N(n8455), .A1N(image_data[112]), 
        .Y(n7540) );
  AOI22XL U6843 ( .A0(n8114), .A1(n8430), .B0(n3384), .B1(n3360), .Y(n7539) );
  AOI211XL U6844 ( .A0(n3351), .A1(n3428), .B0(n7282), .C0(n7281), .Y(n2921)
         );
  AOI2BB2XL U6845 ( .B0(n3346), .B1(n8455), .A0N(n8455), .A1N(image_data[113]), 
        .Y(n7281) );
  AOI22XL U6846 ( .A0(n3384), .A1(n3375), .B0(n8452), .B1(n6332), .Y(n7280) );
  AOI211XL U6847 ( .A0(n7795), .A1(n3428), .B0(n7791), .C0(n7790), .Y(n2922)
         );
  AOI2BB2XL U6848 ( .B0(n3348), .B1(n8455), .A0N(n8455), .A1N(image_data[114]), 
        .Y(n7790) );
  AOI22XL U6849 ( .A0(n8452), .A1(n6880), .B0(n3384), .B1(n3395), .Y(n7789) );
  AOI211XL U6850 ( .A0(n3369), .A1(n3428), .B0(n8457), .C0(n8456), .Y(n2923)
         );
  AOI2BB2XL U6851 ( .B0(n3347), .B1(n8455), .A0N(n8455), .A1N(image_data[115]), 
        .Y(n8456) );
  AOI22XL U6852 ( .A0(n8452), .A1(n6291), .B0(n3384), .B1(n3349), .Y(n8453) );
  AOI211XL U6853 ( .A0(n8503), .A1(n3428), .B0(n7538), .C0(n7537), .Y(n2924)
         );
  AOI2BB2XL U6854 ( .B0(n6855), .B1(n8455), .A0N(n8455), .A1N(image_data[116]), 
        .Y(n7537) );
  AOI22XL U6855 ( .A0(n3371), .A1(n8430), .B0(n3384), .B1(n3388), .Y(n7536) );
  AOI211XL U6856 ( .A0(n3361), .A1(n3428), .B0(n7285), .C0(n7284), .Y(n2925)
         );
  AOI2BB2XL U6857 ( .B0(n8496), .B1(n8455), .A0N(n8455), .A1N(image_data[117]), 
        .Y(n7284) );
  AOI22XL U6858 ( .A0(n3384), .A1(n6979), .B0(n8452), .B1(n7078), .Y(n7283) );
  AOI211XL U6859 ( .A0(n3352), .A1(n3428), .B0(n7622), .C0(n7621), .Y(n2926)
         );
  AOI2BB2XL U6860 ( .B0(n3365), .B1(n8455), .A0N(n8455), .A1N(image_data[118]), 
        .Y(n7621) );
  AOI22XL U6861 ( .A0(n8430), .A1(n3353), .B0(n3384), .B1(n7581), .Y(n7619) );
  AOI211XL U6862 ( .A0(n3362), .A1(n3428), .B0(n6772), .C0(n6771), .Y(n2927)
         );
  AOI2BB2XL U6863 ( .B0(n6586), .B1(n8455), .A0N(n8455), .A1N(image_data[119]), 
        .Y(n6771) );
  AOI22XL U6864 ( .A0(n8452), .A1(n6651), .B0(n3384), .B1(n3368), .Y(n6769) );
  AOI211XL U6865 ( .A0(n3355), .A1(n8397), .B0(n7344), .C0(n7343), .Y(n2928)
         );
  AOI2BB2XL U6866 ( .B0(n3344), .B1(n8394), .A0N(n8394), .A1N(image_data[120]), 
        .Y(n7343) );
  AOI22XL U6867 ( .A0(n6145), .A1(n8452), .B0(n3382), .B1(n3360), .Y(n7342) );
  AOI211XL U6868 ( .A0(n3351), .A1(n8397), .B0(n7115), .C0(n7114), .Y(n2929)
         );
  AOI2BB2XL U6869 ( .B0(n3346), .B1(n8394), .A0N(n8394), .A1N(image_data[121]), 
        .Y(n7114) );
  AOI22XL U6870 ( .A0(n7298), .A1(n8452), .B0(n3382), .B1(n3375), .Y(n7113) );
  AOI211XL U6871 ( .A0(n7795), .A1(n8397), .B0(n7810), .C0(n7809), .Y(n2930)
         );
  AOI2BB2XL U6872 ( .B0(n3348), .B1(n8394), .A0N(n8394), .A1N(image_data[122]), 
        .Y(n7809) );
  AOI22XL U6873 ( .A0(n3358), .A1(n8452), .B0(n3382), .B1(n3395), .Y(n7808) );
  AOI211XL U6874 ( .A0(n3369), .A1(n8397), .B0(n8396), .C0(n8395), .Y(n2931)
         );
  AOI2BB2XL U6875 ( .B0(n3347), .B1(n8394), .A0N(n8394), .A1N(image_data[123]), 
        .Y(n8395) );
  AOI22XL U6876 ( .A0(n8423), .A1(n8452), .B0(n3382), .B1(n3349), .Y(n8392) );
  AOI22XL U6877 ( .A0(n3371), .A1(n8452), .B0(n3382), .B1(n3388), .Y(n5802) );
  AOI211XL U6878 ( .A0(n3361), .A1(n8397), .B0(n7106), .C0(n7105), .Y(n2933)
         );
  AOI2BB2XL U6879 ( .B0(n8496), .B1(n8394), .A0N(n8394), .A1N(image_data[125]), 
        .Y(n7105) );
  AOI22XL U6880 ( .A0(n3357), .A1(n8452), .B0(n3382), .B1(n6979), .Y(n7104) );
  AOI211XL U6881 ( .A0(n3352), .A1(n8397), .B0(n7594), .C0(n7593), .Y(n2934)
         );
  AOI2BB2XL U6882 ( .B0(n3365), .B1(n8394), .A0N(n8394), .A1N(image_data[126]), 
        .Y(n7593) );
  AOI22XL U6883 ( .A0(n8452), .A1(n3353), .B0(n3382), .B1(n7581), .Y(n7592) );
  AOI211XL U6884 ( .A0(n3362), .A1(n8397), .B0(n6613), .C0(n6612), .Y(n2935)
         );
  AOI2BB2XL U6885 ( .B0(n6586), .B1(n8394), .A0N(n8394), .A1N(image_data[127]), 
        .Y(n6612) );
  AOI22XL U6886 ( .A0(n3354), .A1(n8452), .B0(n3382), .B1(n3368), .Y(n6611) );
  AOI211XL U6887 ( .A0(n3355), .A1(n8206), .B0(n7398), .C0(n7397), .Y(n2936)
         );
  AOI2BB2XL U6888 ( .B0(n3344), .B1(n8203), .A0N(n8203), .A1N(image_data[128]), 
        .Y(n7397) );
  AOI22XL U6889 ( .A0(n8200), .A1(n8114), .B0(n8260), .B1(n3356), .Y(n7396) );
  AOI211XL U6890 ( .A0(n3351), .A1(n8206), .B0(n7145), .C0(n7144), .Y(n2937)
         );
  AOI2BB2XL U6891 ( .B0(n3346), .B1(n8203), .A0N(n8203), .A1N(image_data[129]), 
        .Y(n7144) );
  AOI22XL U6892 ( .A0(n7298), .A1(n8200), .B0(n8273), .B1(n3375), .Y(n7143) );
  AOI211XL U6893 ( .A0(n7795), .A1(n8206), .B0(n7825), .C0(n7824), .Y(n2938)
         );
  AOI2BB2XL U6894 ( .B0(n3348), .B1(n8203), .A0N(n8203), .A1N(image_data[130]), 
        .Y(n7824) );
  AOI22XL U6895 ( .A0(n8260), .A1(n6880), .B0(n8273), .B1(n3395), .Y(n7823) );
  AOI211XL U6896 ( .A0(n3369), .A1(n8206), .B0(n8205), .C0(n8204), .Y(n2939)
         );
  AOI2BB2XL U6897 ( .B0(n3347), .B1(n8203), .A0N(n8203), .A1N(image_data[131]), 
        .Y(n8204) );
  AOI22XL U6898 ( .A0(n8423), .A1(n8200), .B0(n8260), .B1(n6291), .Y(n8201) );
  AOI211XL U6899 ( .A0(n8503), .A1(n8206), .B0(n7392), .C0(n7391), .Y(n2940)
         );
  AOI2BB2XL U6900 ( .B0(n6855), .B1(n8203), .A0N(n8203), .A1N(image_data[132]), 
        .Y(n7391) );
  AOI22XL U6901 ( .A0(n3371), .A1(n8200), .B0(n8260), .B1(n7326), .Y(n7390) );
  AOI211XL U6902 ( .A0(n3361), .A1(n8206), .B0(n7139), .C0(n7138), .Y(n2941)
         );
  AOI2BB2XL U6903 ( .B0(n8496), .B1(n8203), .A0N(n8203), .A1N(image_data[133]), 
        .Y(n7138) );
  AOI22XL U6904 ( .A0(n3357), .A1(n8200), .B0(n8273), .B1(n6979), .Y(n7137) );
  AOI211XL U6905 ( .A0(n3352), .A1(n8206), .B0(n7664), .C0(n7663), .Y(n2942)
         );
  AOI2BB2XL U6906 ( .B0(n3365), .B1(n8203), .A0N(n8203), .A1N(image_data[134]), 
        .Y(n7663) );
  AOI22XL U6907 ( .A0(n8273), .A1(n7581), .B0(n8260), .B1(n3350), .Y(n7662) );
  AOI211XL U6908 ( .A0(n3362), .A1(n8206), .B0(n6671), .C0(n6670), .Y(n2943)
         );
  AOI2BB2XL U6909 ( .B0(n6586), .B1(n8203), .A0N(n8203), .A1N(image_data[135]), 
        .Y(n6670) );
  AOI22XL U6910 ( .A0(n8260), .A1(n6651), .B0(n8273), .B1(n3368), .Y(n6669) );
  AOI211XL U6911 ( .A0(n3355), .A1(n8265), .B0(n7434), .C0(n7433), .Y(n2944)
         );
  AOI2BB2XL U6912 ( .B0(n3344), .B1(n8262), .A0N(n8262), .A1N(image_data[136]), 
        .Y(n7433) );
  AOI22XL U6913 ( .A0(n8114), .A1(n8260), .B0(n8141), .B1(n3360), .Y(n7432) );
  AOI211XL U6914 ( .A0(n3351), .A1(n8265), .B0(n7184), .C0(n7183), .Y(n2945)
         );
  AOI2BB2XL U6915 ( .B0(n3366), .B1(n8262), .A0N(n8262), .A1N(image_data[137]), 
        .Y(n7183) );
  AOI22XL U6916 ( .A0(n7298), .A1(n8260), .B0(n8141), .B1(n3375), .Y(n7182) );
  AOI211XL U6917 ( .A0(n7795), .A1(n8265), .B0(n7859), .C0(n7858), .Y(n2946)
         );
  AOI2BB2XL U6918 ( .B0(n3348), .B1(n8262), .A0N(n8262), .A1N(image_data[138]), 
        .Y(n7858) );
  AOI22XL U6919 ( .A0(n3358), .A1(n8260), .B0(n8141), .B1(n3395), .Y(n7857) );
  AOI211XL U6920 ( .A0(n3369), .A1(n8265), .B0(n8264), .C0(n8263), .Y(n2947)
         );
  AOI2BB2XL U6921 ( .B0(n3347), .B1(n8262), .A0N(n8262), .A1N(image_data[139]), 
        .Y(n8263) );
  AOI22XL U6922 ( .A0(n8423), .A1(n8260), .B0(n8259), .B1(n6291), .Y(n8261) );
  AOI211XL U6923 ( .A0(n8503), .A1(n8265), .B0(n7431), .C0(n7430), .Y(n2948)
         );
  AOI2BB2XL U6924 ( .B0(n6855), .B1(n8262), .A0N(n8262), .A1N(image_data[140]), 
        .Y(n7430) );
  AOI22XL U6925 ( .A0(n8141), .A1(n3388), .B0(n8259), .B1(n7326), .Y(n7429) );
  AOI21XL U6926 ( .A0(n3357), .A1(n8260), .B0(n6340), .Y(n2949) );
  AOI2BB2XL U6927 ( .B0(n6339), .B1(n8262), .A0N(n8262), .A1N(image_data[141]), 
        .Y(n6340) );
  OAI22XL U6928 ( .A0(n7963), .A1(n8275), .B0(n7307), .B1(n6682), .Y(n6336) );
  AOI211XL U6929 ( .A0(n3352), .A1(n8265), .B0(n7686), .C0(n7685), .Y(n2950)
         );
  AOI2BB2XL U6930 ( .B0(n3345), .B1(n8262), .A0N(n8262), .A1N(image_data[142]), 
        .Y(n7685) );
  AOI22XL U6931 ( .A0(n8141), .A1(n7581), .B0(n8259), .B1(n3350), .Y(n7683) );
  AOI211XL U6932 ( .A0(n3362), .A1(n8265), .B0(n6686), .C0(n6685), .Y(n2951)
         );
  AOI2BB2XL U6933 ( .B0(n6959), .B1(n8262), .A0N(n8262), .A1N(image_data[143]), 
        .Y(n6685) );
  AOI22XL U6934 ( .A0(n8259), .A1(n6651), .B0(n8141), .B1(n3368), .Y(n6684) );
  AOI211XL U6935 ( .A0(n3355), .A1(n8198), .B0(n7404), .C0(n7403), .Y(n2952)
         );
  AOI2BB2XL U6936 ( .B0(n3344), .B1(n8195), .A0N(n8195), .A1N(image_data[144]), 
        .Y(n7403) );
  AOI22XL U6937 ( .A0(n6145), .A1(n8259), .B0(n3383), .B1(n3360), .Y(n7402) );
  AOI211XL U6938 ( .A0(n3351), .A1(n8198), .B0(n7133), .C0(n7132), .Y(n2953)
         );
  AOI2BB2XL U6939 ( .B0(n3366), .B1(n8195), .A0N(n8195), .A1N(image_data[145]), 
        .Y(n7132) );
  AOI22XL U6940 ( .A0(n7298), .A1(n8259), .B0(n3383), .B1(n3375), .Y(n7131) );
  AOI211XL U6941 ( .A0(n7795), .A1(n8198), .B0(n7838), .C0(n7837), .Y(n2954)
         );
  AOI2BB2XL U6942 ( .B0(n3348), .B1(n8195), .A0N(n8195), .A1N(image_data[146]), 
        .Y(n7837) );
  AOI22XL U6943 ( .A0(n3358), .A1(n8259), .B0(n3383), .B1(n3395), .Y(n7836) );
  AOI211XL U6944 ( .A0(n3369), .A1(n8198), .B0(n8197), .C0(n8196), .Y(n2955)
         );
  AOI2BB2XL U6945 ( .B0(n3347), .B1(n8195), .A0N(n8195), .A1N(image_data[147]), 
        .Y(n8196) );
  AOI22XL U6946 ( .A0(n8404), .A1(n6291), .B0(n3383), .B1(n3349), .Y(n8194) );
  AOI211XL U6947 ( .A0(n8503), .A1(n8198), .B0(n7380), .C0(n7379), .Y(n2956)
         );
  AOI2BB2XL U6948 ( .B0(n6855), .B1(n8195), .A0N(n8195), .A1N(image_data[148]), 
        .Y(n7379) );
  AOI22XL U6949 ( .A0(n3383), .A1(n3388), .B0(n8404), .B1(n7326), .Y(n7378) );
  AOI211XL U6950 ( .A0(n3361), .A1(n8198), .B0(n7130), .C0(n7129), .Y(n2957)
         );
  AOI2BB2XL U6951 ( .B0(n8496), .B1(n8195), .A0N(n8195), .A1N(image_data[149]), 
        .Y(n7129) );
  AOI22XL U6952 ( .A0(n3357), .A1(n8259), .B0(n3383), .B1(n6979), .Y(n7128) );
  AOI211XL U6953 ( .A0(n3352), .A1(n8198), .B0(n7655), .C0(n7654), .Y(n2958)
         );
  AOI2BB2XL U6954 ( .B0(n3365), .B1(n8195), .A0N(n8195), .A1N(image_data[150]), 
        .Y(n7654) );
  AOI22XL U6955 ( .A0(n8259), .A1(n3353), .B0(n3383), .B1(n7581), .Y(n7653) );
  AOI211XL U6956 ( .A0(n3362), .A1(n8198), .B0(n6619), .C0(n6618), .Y(n2959)
         );
  AOI2BB2XL U6957 ( .B0(n6586), .B1(n8195), .A0N(n8195), .A1N(image_data[151]), 
        .Y(n6618) );
  AOI22XL U6958 ( .A0(n3354), .A1(n8259), .B0(n3383), .B1(n3368), .Y(n6617) );
  AOI211XL U6959 ( .A0(n3355), .A1(n8213), .B0(n7407), .C0(n7406), .Y(n2960)
         );
  AOI2BB2XL U6960 ( .B0(n3344), .B1(n8210), .A0N(n8210), .A1N(image_data[152]), 
        .Y(n7406) );
  AOI22XL U6961 ( .A0(n8114), .A1(n8404), .B0(n3377), .B1(n3360), .Y(n7405) );
  AOI211XL U6962 ( .A0(n3351), .A1(n8213), .B0(n7148), .C0(n7147), .Y(n2961)
         );
  AOI2BB2XL U6963 ( .B0(n3346), .B1(n8210), .A0N(n8210), .A1N(image_data[153]), 
        .Y(n7147) );
  AOI22XL U6964 ( .A0(n7298), .A1(n8404), .B0(n3377), .B1(n3375), .Y(n7146) );
  AOI211XL U6965 ( .A0(n7795), .A1(n8213), .B0(n7835), .C0(n7834), .Y(n2962)
         );
  AOI2BB2XL U6966 ( .B0(n3348), .B1(n8210), .A0N(n8210), .A1N(image_data[154]), 
        .Y(n7834) );
  AOI22XL U6967 ( .A0(n3358), .A1(n8404), .B0(n3377), .B1(n3395), .Y(n7833) );
  AOI211XL U6968 ( .A0(n3369), .A1(n8213), .B0(n8212), .C0(n8211), .Y(n2963)
         );
  AOI2BB2XL U6969 ( .B0(n3347), .B1(n8210), .A0N(n8210), .A1N(image_data[155]), 
        .Y(n8211) );
  AOI22XL U6970 ( .A0(n8207), .A1(n6291), .B0(n3377), .B1(n3349), .Y(n8208) );
  AOI211XL U6971 ( .A0(n8503), .A1(n8213), .B0(n7376), .C0(n7375), .Y(n2964)
         );
  AOI2BB2XL U6972 ( .B0(n6855), .B1(n8210), .A0N(n8210), .A1N(image_data[156]), 
        .Y(n7375) );
  AOI22XL U6973 ( .A0(n3371), .A1(n8404), .B0(n3377), .B1(n3388), .Y(n7374) );
  AOI211XL U6974 ( .A0(n3361), .A1(n8213), .B0(n7124), .C0(n7123), .Y(n2965)
         );
  AOI2BB2XL U6975 ( .B0(n8496), .B1(n8210), .A0N(n8210), .A1N(image_data[157]), 
        .Y(n7123) );
  AOI22XL U6976 ( .A0(n3377), .A1(n6979), .B0(n8207), .B1(n7078), .Y(n7122) );
  AOI211XL U6977 ( .A0(n3352), .A1(n8213), .B0(n7649), .C0(n7648), .Y(n2966)
         );
  AOI2BB2XL U6978 ( .B0(n3345), .B1(n8210), .A0N(n8210), .A1N(image_data[158]), 
        .Y(n7648) );
  AOI22XL U6979 ( .A0(n3377), .A1(n7581), .B0(n8207), .B1(n3350), .Y(n7647) );
  AOI211XL U6980 ( .A0(n3362), .A1(n8213), .B0(n6630), .C0(n6629), .Y(n2967)
         );
  AOI2BB2XL U6981 ( .B0(n6959), .B1(n8210), .A0N(n8210), .A1N(image_data[159]), 
        .Y(n6629) );
  AOI22XL U6982 ( .A0(n3354), .A1(n8404), .B0(n3377), .B1(n3368), .Y(n6628) );
  AOI211XL U6983 ( .A0(n3355), .A1(n3427), .B0(n7478), .C0(n7477), .Y(n2968)
         );
  AOI2BB2XL U6984 ( .B0(n3344), .B1(n8305), .A0N(n8305), .A1N(image_data[160]), 
        .Y(n7477) );
  AOI22XL U6985 ( .A0(n8114), .A1(n8207), .B0(n8301), .B1(n3360), .Y(n7476) );
  AOI211XL U6986 ( .A0(n3351), .A1(n3427), .B0(n7236), .C0(n7235), .Y(n2969)
         );
  AOI2BB2XL U6987 ( .B0(n3346), .B1(n8305), .A0N(n8305), .A1N(image_data[161]), 
        .Y(n7235) );
  AOI22XL U6988 ( .A0(n7298), .A1(n8207), .B0(n8301), .B1(n3375), .Y(n7234) );
  AOI211XL U6989 ( .A0(n7795), .A1(n3427), .B0(n7872), .C0(n7871), .Y(n2970)
         );
  AOI2BB2XL U6990 ( .B0(n3348), .B1(n8305), .A0N(n8305), .A1N(image_data[162]), 
        .Y(n7871) );
  AOI22XL U6991 ( .A0(n7923), .A1(n8207), .B0(n8301), .B1(n3395), .Y(n7870) );
  AOI211XL U6992 ( .A0(n3369), .A1(n3427), .B0(n8307), .C0(n8306), .Y(n2971)
         );
  AOI2BB2XL U6993 ( .B0(n3347), .B1(n8305), .A0N(n8305), .A1N(image_data[163]), 
        .Y(n8306) );
  AOI22XL U6994 ( .A0(n8302), .A1(n6291), .B0(n8301), .B1(n3349), .Y(n8303) );
  AOI211XL U6995 ( .A0(n8503), .A1(n3427), .B0(n7481), .C0(n7480), .Y(n2972)
         );
  AOI2BB2XL U6996 ( .B0(n6855), .B1(n8305), .A0N(n8305), .A1N(image_data[164]), 
        .Y(n7480) );
  AOI22XL U6997 ( .A0(n3371), .A1(n8207), .B0(n8301), .B1(n3388), .Y(n7479) );
  AOI211XL U6998 ( .A0(n3361), .A1(n3427), .B0(n7230), .C0(n7229), .Y(n2973)
         );
  AOI2BB2XL U6999 ( .B0(n8496), .B1(n8305), .A0N(n8305), .A1N(image_data[165]), 
        .Y(n7229) );
  AOI22XL U7000 ( .A0(n3357), .A1(n8207), .B0(n8301), .B1(n6979), .Y(n7228) );
  AOI211XL U7001 ( .A0(n3352), .A1(n3427), .B0(n7704), .C0(n7703), .Y(n2974)
         );
  AOI2BB2XL U7002 ( .B0(n3345), .B1(n8305), .A0N(n8305), .A1N(image_data[166]), 
        .Y(n7703) );
  AOI22XL U7003 ( .A0(n8207), .A1(n3353), .B0(n8302), .B1(n3350), .Y(n7702) );
  AOI211XL U7004 ( .A0(n3362), .A1(n3427), .B0(n6725), .C0(n6724), .Y(n2975)
         );
  AOI2BB2XL U7005 ( .B0(n6586), .B1(n8305), .A0N(n8305), .A1N(image_data[167]), 
        .Y(n6724) );
  AOI22XL U7006 ( .A0(n3354), .A1(n8207), .B0(n8301), .B1(n3368), .Y(n6722) );
  AOI211XL U7007 ( .A0(n3355), .A1(n8367), .B0(n7544), .C0(n7543), .Y(n2976)
         );
  AOI2BB2XL U7008 ( .B0(n3344), .B1(n8364), .A0N(n8364), .A1N(image_data[168]), 
        .Y(n7543) );
  AOI22XL U7009 ( .A0(n8362), .A1(n3360), .B0(n3384), .B1(n3356), .Y(n7542) );
  AOI211XL U7010 ( .A0(n3351), .A1(n8367), .B0(n7288), .C0(n7287), .Y(n2977)
         );
  AOI2BB2XL U7011 ( .B0(n3366), .B1(n8364), .A0N(n8364), .A1N(image_data[169]), 
        .Y(n7287) );
  AOI22XL U7012 ( .A0(n8362), .A1(n3375), .B0(n3384), .B1(n6332), .Y(n7286) );
  AOI211XL U7013 ( .A0(n7795), .A1(n8367), .B0(n7916), .C0(n7915), .Y(n2978)
         );
  AOI2BB2XL U7014 ( .B0(n3348), .B1(n8364), .A0N(n8364), .A1N(image_data[170]), 
        .Y(n7915) );
  AOI22XL U7015 ( .A0(n3384), .A1(n6880), .B0(n8362), .B1(n3395), .Y(n7914) );
  AOI211XL U7016 ( .A0(n3369), .A1(n8367), .B0(n8366), .C0(n8365), .Y(n2979)
         );
  AOI2BB2XL U7017 ( .B0(n3347), .B1(n8364), .A0N(n8364), .A1N(image_data[171]), 
        .Y(n8365) );
  AOI22XL U7018 ( .A0(n3384), .A1(n6291), .B0(n8362), .B1(n3349), .Y(n8363) );
  AOI211XL U7019 ( .A0(n8503), .A1(n8367), .B0(n7553), .C0(n7552), .Y(n2980)
         );
  AOI2BB2XL U7020 ( .B0(n6855), .B1(n8364), .A0N(n8364), .A1N(image_data[172]), 
        .Y(n7552) );
  AOI22XL U7021 ( .A0(n8362), .A1(n3388), .B0(n3384), .B1(n7326), .Y(n7551) );
  AOI211XL U7022 ( .A0(n3361), .A1(n8367), .B0(n7294), .C0(n7293), .Y(n2981)
         );
  AOI2BB2XL U7023 ( .B0(n8496), .B1(n8364), .A0N(n8364), .A1N(image_data[173]), 
        .Y(n7293) );
  AOI22XL U7024 ( .A0(n8362), .A1(n6979), .B0(n3384), .B1(n7078), .Y(n7292) );
  AOI211XL U7025 ( .A0(n3352), .A1(n8367), .B0(n7738), .C0(n7737), .Y(n2982)
         );
  AOI2BB2XL U7026 ( .B0(n3345), .B1(n8364), .A0N(n8364), .A1N(image_data[174]), 
        .Y(n7737) );
  AOI22XL U7027 ( .A0(n8362), .A1(n7581), .B0(n3384), .B1(n3350), .Y(n7736) );
  AOI211XL U7028 ( .A0(n3362), .A1(n8367), .B0(n6784), .C0(n6783), .Y(n2983)
         );
  AOI2BB2XL U7029 ( .B0(n6586), .B1(n8364), .A0N(n8364), .A1N(image_data[175]), 
        .Y(n6783) );
  AOI22XL U7030 ( .A0(n3384), .A1(n6651), .B0(n8362), .B1(n3368), .Y(n6781) );
  AOI211XL U7031 ( .A0(n3355), .A1(n7922), .B0(n7547), .C0(n7546), .Y(n2984)
         );
  AOI2BB2XL U7032 ( .B0(n3344), .B1(n7919), .A0N(n7919), .A1N(image_data[176]), 
        .Y(n7546) );
  AOI22XL U7033 ( .A0(n3384), .A1(n8114), .B0(n3382), .B1(n3356), .Y(n7545) );
  AOI211XL U7034 ( .A0(n3351), .A1(n7922), .B0(n7291), .C0(n7290), .Y(n2985)
         );
  AOI2BB2XL U7035 ( .B0(n3366), .B1(n7919), .A0N(n7919), .A1N(image_data[177]), 
        .Y(n7290) );
  AOI22XL U7036 ( .A0(n3384), .A1(n7298), .B0(n3382), .B1(n6332), .Y(n7289) );
  AOI211XL U7037 ( .A0(n7795), .A1(n7922), .B0(n7921), .C0(n7920), .Y(n2986)
         );
  AOI2BB2XL U7038 ( .B0(n3348), .B1(n7919), .A0N(n7919), .A1N(image_data[178]), 
        .Y(n7920) );
  AOI22XL U7039 ( .A0(n3358), .A1(n3384), .B0(n3382), .B1(n6880), .Y(n7917) );
  AOI22XL U7040 ( .A0(n8423), .A1(n3384), .B0(n3382), .B1(n6291), .Y(n6292) );
  AOI211XL U7041 ( .A0(n8503), .A1(n7922), .B0(n7550), .C0(n7549), .Y(n2988)
         );
  AOI2BB2XL U7042 ( .B0(n6855), .B1(n7919), .A0N(n7919), .A1N(image_data[180]), 
        .Y(n7549) );
  AOI22XL U7043 ( .A0(n3371), .A1(n3384), .B0(n3382), .B1(n7326), .Y(n7548) );
  AOI211XL U7044 ( .A0(n3361), .A1(n7922), .B0(n7297), .C0(n7296), .Y(n2989)
         );
  AOI2BB2XL U7045 ( .B0(n8496), .B1(n7919), .A0N(n7919), .A1N(image_data[181]), 
        .Y(n7296) );
  AOI22XL U7046 ( .A0(n3357), .A1(n3384), .B0(n3382), .B1(n7078), .Y(n7295) );
  AOI211XL U7047 ( .A0(n3352), .A1(n7922), .B0(n7742), .C0(n7741), .Y(n2990)
         );
  AOI2BB2XL U7048 ( .B0(n3365), .B1(n7919), .A0N(n7919), .A1N(image_data[182]), 
        .Y(n7741) );
  AOI22XL U7049 ( .A0(n3384), .A1(n3353), .B0(n3382), .B1(n3350), .Y(n7739) );
  AOI211XL U7050 ( .A0(n3362), .A1(n7922), .B0(n6775), .C0(n6774), .Y(n2991)
         );
  AOI2BB2XL U7051 ( .B0(n6586), .B1(n7919), .A0N(n7919), .A1N(image_data[183]), 
        .Y(n6774) );
  AOI22XL U7052 ( .A0(n3354), .A1(n3384), .B0(n3382), .B1(n6651), .Y(n6773) );
  AOI221XL U7053 ( .A0(image_data[184]), .A1(n7569), .B0(n6990), .B1(n8148), 
        .C0(n6989), .Y(n2992) );
  AOI211XL U7054 ( .A0(n3351), .A1(n8151), .B0(n7074), .C0(n7073), .Y(n2993)
         );
  AOI2BB2XL U7055 ( .B0(n3346), .B1(n8148), .A0N(n8148), .A1N(image_data[185]), 
        .Y(n7073) );
  AOI22XL U7056 ( .A0(n3382), .A1(n7298), .B0(n8273), .B1(n6332), .Y(n7072) );
  AOI211XL U7057 ( .A0(n7795), .A1(n8151), .B0(n7798), .C0(n7797), .Y(n2994)
         );
  AOI2BB2XL U7058 ( .B0(n3348), .B1(n8148), .A0N(n8148), .A1N(image_data[186]), 
        .Y(n7797) );
  AOI22XL U7059 ( .A0(n3358), .A1(n3382), .B0(n8273), .B1(n6880), .Y(n7796) );
  AOI211XL U7060 ( .A0(n3369), .A1(n8151), .B0(n8150), .C0(n8149), .Y(n2995)
         );
  AOI2BB2XL U7061 ( .B0(n3347), .B1(n8148), .A0N(n8148), .A1N(image_data[187]), 
        .Y(n8149) );
  AOI22XL U7062 ( .A0(n8423), .A1(n3382), .B0(n8273), .B1(n6291), .Y(n8147) );
  AOI211XL U7063 ( .A0(n8503), .A1(n8151), .B0(n7329), .C0(n7328), .Y(n2996)
         );
  AOI2BB2XL U7064 ( .B0(n6855), .B1(n8148), .A0N(n8148), .A1N(image_data[188]), 
        .Y(n7328) );
  AOI22XL U7065 ( .A0(n3371), .A1(n3382), .B0(n8273), .B1(n7326), .Y(n7327) );
  AOI211XL U7066 ( .A0(n3361), .A1(n8151), .B0(n7081), .C0(n7080), .Y(n2997)
         );
  AOI2BB2XL U7067 ( .B0(n8496), .B1(n8148), .A0N(n8148), .A1N(image_data[189]), 
        .Y(n7080) );
  AOI22XL U7068 ( .A0(n3357), .A1(n3382), .B0(n8273), .B1(n7078), .Y(n7079) );
  AOI211XL U7069 ( .A0(n3352), .A1(n8151), .B0(n7634), .C0(n7633), .Y(n2998)
         );
  AOI2BB2XL U7070 ( .B0(n3345), .B1(n8148), .A0N(n8148), .A1N(image_data[190]), 
        .Y(n7633) );
  AOI22XL U7071 ( .A0(n3382), .A1(n3353), .B0(n8273), .B1(n3350), .Y(n7632) );
  AOI221XL U7072 ( .A0(image_data[191]), .A1(n7569), .B0(n7568), .B1(n8148), 
        .C0(n7567), .Y(n2999) );
  AOI22XL U7073 ( .A0(n3354), .A1(n3382), .B0(n8273), .B1(n6651), .Y(n7565) );
  AOI211XL U7074 ( .A0(n3355), .A1(n8279), .B0(n7447), .C0(n7446), .Y(n3000)
         );
  AOI2BB2XL U7075 ( .B0(n3344), .B1(n8276), .A0N(n8276), .A1N(image_data[192]), 
        .Y(n7446) );
  AOI22XL U7076 ( .A0(n8114), .A1(n8273), .B0(n3378), .B1(n3360), .Y(n7444) );
  AOI211XL U7077 ( .A0(n3351), .A1(n8279), .B0(n7206), .C0(n7205), .Y(n3001)
         );
  AOI2BB2XL U7078 ( .B0(n3346), .B1(n8276), .A0N(n8276), .A1N(image_data[193]), 
        .Y(n7205) );
  AOI22XL U7079 ( .A0(n7298), .A1(n8273), .B0(n3378), .B1(n3375), .Y(n7204) );
  AOI211XL U7080 ( .A0(n7795), .A1(n8279), .B0(n7862), .C0(n7861), .Y(n3002)
         );
  AOI2BB2XL U7081 ( .B0(n3348), .B1(n8276), .A0N(n8276), .A1N(image_data[194]), 
        .Y(n7861) );
  AOI22XL U7082 ( .A0(n3358), .A1(n8273), .B0(n3378), .B1(n3395), .Y(n7860) );
  AOI211XL U7083 ( .A0(n3369), .A1(n8279), .B0(n8278), .C0(n8277), .Y(n3003)
         );
  AOI2BB2XL U7084 ( .B0(n3347), .B1(n8276), .A0N(n8276), .A1N(image_data[195]), 
        .Y(n8277) );
  AOI22XL U7085 ( .A0(n8423), .A1(n8273), .B0(n3378), .B1(n3349), .Y(n8274) );
  AOI211XL U7086 ( .A0(n8503), .A1(n8279), .B0(n7450), .C0(n7449), .Y(n3004)
         );
  AOI2BB2XL U7087 ( .B0(n6855), .B1(n8276), .A0N(n8276), .A1N(image_data[196]), 
        .Y(n7449) );
  AOI22XL U7088 ( .A0(n3371), .A1(n8273), .B0(n3378), .B1(n3388), .Y(n7448) );
  AOI211XL U7089 ( .A0(n3361), .A1(n8279), .B0(n7203), .C0(n7202), .Y(n3005)
         );
  AOI2BB2XL U7090 ( .B0(n8496), .B1(n8276), .A0N(n8276), .A1N(image_data[197]), 
        .Y(n7202) );
  AOI22XL U7091 ( .A0(n3357), .A1(n8273), .B0(n3378), .B1(n6979), .Y(n7201) );
  AOI211XL U7092 ( .A0(n3352), .A1(n8279), .B0(n7689), .C0(n7688), .Y(n3006)
         );
  AOI2BB2XL U7093 ( .B0(n3365), .B1(n8276), .A0N(n8276), .A1N(image_data[198]), 
        .Y(n7688) );
  AOI22XL U7094 ( .A0(n8273), .A1(n3353), .B0(n3378), .B1(n7581), .Y(n7687) );
  AOI211XL U7095 ( .A0(n3362), .A1(n8279), .B0(n6693), .C0(n6692), .Y(n3007)
         );
  AOI2BB2XL U7096 ( .B0(n6586), .B1(n8276), .A0N(n8276), .A1N(image_data[199]), 
        .Y(n6692) );
  AOI22XL U7097 ( .A0(n3354), .A1(n8273), .B0(n3378), .B1(n6787), .Y(n6690) );
  AOI21XL U7098 ( .A0(n3373), .A1(n8146), .B0(n6149), .Y(n3008) );
  AOI22XL U7099 ( .A0(n7898), .A1(n3360), .B0(n3383), .B1(n3356), .Y(n6147) );
  AOI211XL U7100 ( .A0(n7987), .A1(image_data[201]), .B0(n7986), .C0(n7985), 
        .Y(n3009) );
  OAI22XL U7101 ( .A0(n3359), .A1(n8351), .B0(n3374), .B1(n8275), .Y(n7985) );
  AOI21XL U7102 ( .A0(n3366), .A1(n7984), .B0(n7987), .Y(n7986) );
  AOI22XL U7103 ( .A0(n3351), .A1(n7983), .B0(n3383), .B1(n6332), .Y(n7984) );
  AOI211XL U7104 ( .A0(n7795), .A1(n8146), .B0(n7801), .C0(n7800), .Y(n3010)
         );
  AOI2BB2XL U7105 ( .B0(n3348), .B1(n8143), .A0N(n8143), .A1N(image_data[202]), 
        .Y(n7800) );
  AOI22XL U7106 ( .A0(n3358), .A1(n8141), .B0(n3383), .B1(n6880), .Y(n7799) );
  AOI211XL U7107 ( .A0(n3369), .A1(n8146), .B0(n8145), .C0(n8144), .Y(n3011)
         );
  AOI2BB2XL U7108 ( .B0(n3347), .B1(n8143), .A0N(n8143), .A1N(image_data[203]), 
        .Y(n8144) );
  AOI22XL U7109 ( .A0(n8423), .A1(n8141), .B0(n3383), .B1(n6291), .Y(n8142) );
  AOI211XL U7110 ( .A0(n8503), .A1(n8146), .B0(n7332), .C0(n7331), .Y(n3012)
         );
  AOI2BB2XL U7111 ( .B0(n6855), .B1(n8143), .A0N(n8143), .A1N(image_data[204]), 
        .Y(n7331) );
  AOI22XL U7112 ( .A0(n3371), .A1(n8141), .B0(n3383), .B1(n7326), .Y(n7330) );
  AOI211XL U7113 ( .A0(n3361), .A1(n8146), .B0(n7084), .C0(n7083), .Y(n3013)
         );
  AOI2BB2XL U7114 ( .B0(n7303), .B1(n8143), .A0N(n8143), .A1N(image_data[205]), 
        .Y(n7083) );
  AOI22XL U7115 ( .A0(n3357), .A1(n8141), .B0(n3383), .B1(n7078), .Y(n7082) );
  AOI211XL U7116 ( .A0(n3352), .A1(n8146), .B0(n7637), .C0(n7636), .Y(n3014)
         );
  AOI2BB2XL U7117 ( .B0(n3365), .B1(n8143), .A0N(n8143), .A1N(image_data[206]), 
        .Y(n7636) );
  AOI22XL U7118 ( .A0(n8141), .A1(n3353), .B0(n3383), .B1(n3350), .Y(n7635) );
  AOI211XL U7119 ( .A0(n3362), .A1(n8146), .B0(n6591), .C0(n6590), .Y(n3015)
         );
  AOI2BB2XL U7120 ( .B0(n6959), .B1(n8143), .A0N(n8143), .A1N(image_data[207]), 
        .Y(n6590) );
  AOI22XL U7121 ( .A0(n3354), .A1(n8141), .B0(n3383), .B1(n6651), .Y(n6589) );
  AOI211XL U7122 ( .A0(n3355), .A1(n8175), .B0(n7338), .C0(n7337), .Y(n3016)
         );
  AOI2BB2XL U7123 ( .B0(n3344), .B1(n8172), .A0N(n8172), .A1N(image_data[208]), 
        .Y(n7337) );
  AOI22XL U7124 ( .A0(n3383), .A1(n8114), .B0(n3377), .B1(n3356), .Y(n7336) );
  AOI211XL U7125 ( .A0(n3351), .A1(n8175), .B0(n7112), .C0(n7111), .Y(n3017)
         );
  AOI2BB2XL U7126 ( .B0(n3346), .B1(n8172), .A0N(n8172), .A1N(image_data[209]), 
        .Y(n7111) );
  AOI22XL U7127 ( .A0(n3383), .A1(n7298), .B0(n3377), .B1(n6332), .Y(n7110) );
  AOI211XL U7128 ( .A0(n7795), .A1(n8175), .B0(n7816), .C0(n7815), .Y(n3018)
         );
  AOI2BB2XL U7129 ( .B0(n3348), .B1(n8172), .A0N(n8172), .A1N(image_data[210]), 
        .Y(n7815) );
  AOI22XL U7130 ( .A0(n3358), .A1(n3383), .B0(n3377), .B1(n6880), .Y(n7814) );
  AOI211XL U7131 ( .A0(n3369), .A1(n8175), .B0(n8174), .C0(n8173), .Y(n3019)
         );
  AOI2BB2XL U7132 ( .B0(n3347), .B1(n8172), .A0N(n8172), .A1N(image_data[211]), 
        .Y(n8173) );
  AOI22XL U7133 ( .A0(n8423), .A1(n3383), .B0(n3377), .B1(n6291), .Y(n8170) );
  AOI211XL U7134 ( .A0(n8503), .A1(n8175), .B0(n7364), .C0(n7363), .Y(n3020)
         );
  AOI2BB2XL U7135 ( .B0(n6855), .B1(n8172), .A0N(n8172), .A1N(image_data[212]), 
        .Y(n7363) );
  AOI22XL U7136 ( .A0(n3371), .A1(n3383), .B0(n3377), .B1(n7326), .Y(n7362) );
  AOI211XL U7137 ( .A0(n3361), .A1(n8175), .B0(n7118), .C0(n7117), .Y(n3021)
         );
  AOI2BB2XL U7138 ( .B0(n7303), .B1(n8172), .A0N(n8172), .A1N(image_data[213]), 
        .Y(n7117) );
  AOI22XL U7139 ( .A0(n3357), .A1(n3383), .B0(n3377), .B1(n7078), .Y(n7116) );
  AOI21XL U7140 ( .A0(n3352), .A1(n8175), .B0(n6164), .Y(n3022) );
  AOI22XL U7141 ( .A0(n6143), .A1(n7581), .B0(n3377), .B1(n3350), .Y(n6161) );
  AOI211XL U7142 ( .A0(n3362), .A1(n8175), .B0(n6604), .C0(n6603), .Y(n3023)
         );
  AOI2BB2XL U7143 ( .B0(n6959), .B1(n8172), .A0N(n8172), .A1N(image_data[215]), 
        .Y(n6603) );
  AOI22XL U7144 ( .A0(n3354), .A1(n3383), .B0(n3377), .B1(n6651), .Y(n6602) );
  AOI211XL U7145 ( .A0(n8181), .A1(n3373), .B0(n6936), .C0(n6935), .Y(n3024)
         );
  NOR2XL U7146 ( .A(n7507), .B(n7907), .Y(n6936) );
  AOI32XL U7147 ( .A0(n3367), .A1(n8178), .A2(n6934), .B0(n6980), .B1(n8555), 
        .Y(n6935) );
  AOI22XL U7148 ( .A0(n3377), .A1(n8114), .B0(n8301), .B1(n3356), .Y(n6934) );
  AOI21XL U7149 ( .A0(n3351), .A1(n8181), .B0(n5927), .Y(n3025) );
  AOI22XL U7150 ( .A0(n3377), .A1(n7298), .B0(n8301), .B1(n6332), .Y(n5925) );
  AOI211XL U7151 ( .A0(n7795), .A1(n8181), .B0(n7813), .C0(n7812), .Y(n3026)
         );
  AOI2BB2XL U7152 ( .B0(n3348), .B1(n8178), .A0N(n8178), .A1N(image_data[218]), 
        .Y(n7812) );
  AOI22XL U7153 ( .A0(n3358), .A1(n3377), .B0(n8501), .B1(n3395), .Y(n7811) );
  AOI211XL U7154 ( .A0(n3369), .A1(n8181), .B0(n8180), .C0(n8179), .Y(n3027)
         );
  AOI2BB2XL U7155 ( .B0(n3347), .B1(n8178), .A0N(n8178), .A1N(image_data[219]), 
        .Y(n8179) );
  AOI22XL U7156 ( .A0(n8423), .A1(n3377), .B0(n8501), .B1(n3349), .Y(n8176) );
  AOI21XL U7157 ( .A0(n8503), .A1(n8181), .B0(n6026), .Y(n3028) );
  AOI22XL U7158 ( .A0(n3371), .A1(n3377), .B0(n8501), .B1(n6852), .Y(n6024) );
  AOI211XL U7159 ( .A0(n8181), .A1(n3361), .B0(n6983), .C0(n6982), .Y(n3029)
         );
  NOR2XL U7160 ( .A(n7956), .B(n8177), .Y(n6983) );
  AOI32XL U7161 ( .A0(n7303), .A1(n8178), .A2(n6981), .B0(n6980), .B1(n8554), 
        .Y(n6982) );
  AOI22XL U7162 ( .A0(n3357), .A1(n3377), .B0(n8501), .B1(n6979), .Y(n6981) );
  AOI211XL U7163 ( .A0(n3352), .A1(n8181), .B0(n7643), .C0(n7642), .Y(n3030)
         );
  AOI2BB2XL U7164 ( .B0(n3345), .B1(n8178), .A0N(n8178), .A1N(image_data[222]), 
        .Y(n7642) );
  AOI22XL U7165 ( .A0(n3377), .A1(n3353), .B0(n8301), .B1(n3350), .Y(n7641) );
  AOI211XL U7166 ( .A0(n3362), .A1(n8181), .B0(n6598), .C0(n6597), .Y(n3031)
         );
  AOI2BB2XL U7167 ( .B0(n6586), .B1(n8178), .A0N(n8178), .A1N(image_data[223]), 
        .Y(n6597) );
  AOI22XL U7168 ( .A0(n3354), .A1(n3377), .B0(n8301), .B1(n6651), .Y(n6596) );
  AOI21XL U7169 ( .A0(n3373), .A1(n8157), .B0(n6141), .Y(n3032) );
  AOI22XL U7170 ( .A0(n8301), .A1(n8114), .B0(n8362), .B1(n3356), .Y(n6139) );
  AOI211XL U7171 ( .A0(n7978), .A1(image_data[225]), .B0(n7977), .C0(n7976), 
        .Y(n3033) );
  OAI22XL U7172 ( .A0(n3359), .A1(n7975), .B0(n3374), .B1(n8177), .Y(n7976) );
  AOI21XL U7173 ( .A0(n3366), .A1(n7974), .B0(n7978), .Y(n7977) );
  AOI22XL U7174 ( .A0(n7973), .A1(n7972), .B0(n8362), .B1(n6332), .Y(n7974) );
  AOI211XL U7175 ( .A0(n7795), .A1(n8157), .B0(n7807), .C0(n7806), .Y(n3034)
         );
  AOI2BB2XL U7176 ( .B0(n3348), .B1(n8154), .A0N(n8154), .A1N(image_data[226]), 
        .Y(n7806) );
  AOI22XL U7177 ( .A0(n3358), .A1(n8301), .B0(n8499), .B1(n3395), .Y(n7805) );
  AOI211XL U7178 ( .A0(n3369), .A1(n8157), .B0(n8156), .C0(n8155), .Y(n3035)
         );
  AOI2BB2XL U7179 ( .B0(n3347), .B1(n8154), .A0N(n8154), .A1N(image_data[227]), 
        .Y(n8155) );
  AOI22XL U7180 ( .A0(n3389), .A1(n8301), .B0(n8499), .B1(n3349), .Y(n8152) );
  AOI211XL U7181 ( .A0(n8503), .A1(n8157), .B0(n7335), .C0(n7334), .Y(n3036)
         );
  AOI2BB2XL U7182 ( .B0(n6855), .B1(n8154), .A0N(n8154), .A1N(image_data[228]), 
        .Y(n7334) );
  AOI22XL U7183 ( .A0(n3371), .A1(n8301), .B0(n8499), .B1(n6852), .Y(n7333) );
  AOI211XL U7184 ( .A0(n3361), .A1(n8157), .B0(n7077), .C0(n7076), .Y(n3037)
         );
  AOI2BB2XL U7185 ( .B0(n7303), .B1(n8154), .A0N(n8154), .A1N(image_data[229]), 
        .Y(n7076) );
  AOI22XL U7186 ( .A0(n3357), .A1(n8301), .B0(n8499), .B1(n6979), .Y(n7075) );
  AOI211XL U7187 ( .A0(n3352), .A1(n8157), .B0(n7631), .C0(n7630), .Y(n3038)
         );
  AOI2BB2XL U7188 ( .B0(n3345), .B1(n8154), .A0N(n8154), .A1N(image_data[230]), 
        .Y(n7630) );
  AOI22XL U7189 ( .A0(n8301), .A1(n3353), .B0(n8499), .B1(n7581), .Y(n7629) );
  AOI211XL U7190 ( .A0(n3362), .A1(n8157), .B0(n6588), .C0(n6587), .Y(n3039)
         );
  AOI2BB2XL U7191 ( .B0(n6959), .B1(n8154), .A0N(n8154), .A1N(image_data[231]), 
        .Y(n6587) );
  AOI22XL U7192 ( .A0(n3354), .A1(n8301), .B0(n8499), .B1(n6787), .Y(n6422) );
  AOI211XL U7193 ( .A0(n3355), .A1(n8293), .B0(n7463), .C0(n7462), .Y(n3040)
         );
  AOI2BB2XL U7194 ( .B0(n3344), .B1(n8290), .A0N(n8290), .A1N(image_data[232]), 
        .Y(n7462) );
  AOI22XL U7195 ( .A0(n8362), .A1(n8114), .B0(n8287), .B1(n3356), .Y(n7461) );
  AOI211XL U7196 ( .A0(n3351), .A1(n8293), .B0(n7218), .C0(n7217), .Y(n3041)
         );
  AOI2BB2XL U7197 ( .B0(n3346), .B1(n8290), .A0N(n8290), .A1N(image_data[233]), 
        .Y(n7217) );
  AOI22XL U7198 ( .A0(n8362), .A1(n7298), .B0(n8287), .B1(n6332), .Y(n7216) );
  AOI211XL U7199 ( .A0(n7795), .A1(n8293), .B0(n7869), .C0(n7868), .Y(n3042)
         );
  AOI2BB2XL U7200 ( .B0(n3348), .B1(n8290), .A0N(n8290), .A1N(image_data[234]), 
        .Y(n7868) );
  AOI22XL U7201 ( .A0(n7923), .A1(n8362), .B0(n8287), .B1(n6880), .Y(n7867) );
  AOI211XL U7202 ( .A0(n3369), .A1(n8293), .B0(n8292), .C0(n8291), .Y(n3043)
         );
  AOI2BB2XL U7203 ( .B0(n3347), .B1(n8290), .A0N(n8290), .A1N(image_data[235]), 
        .Y(n8291) );
  AOI22XL U7204 ( .A0(n8423), .A1(n8362), .B0(n8287), .B1(n6291), .Y(n8288) );
  AOI211XL U7205 ( .A0(n8503), .A1(n8293), .B0(n7469), .C0(n7468), .Y(n3044)
         );
  AOI2BB2XL U7206 ( .B0(n6855), .B1(n8290), .A0N(n8290), .A1N(image_data[236]), 
        .Y(n7468) );
  AOI22XL U7207 ( .A0(n3371), .A1(n8362), .B0(n8287), .B1(n7326), .Y(n7467) );
  AOI211XL U7208 ( .A0(n3361), .A1(n8293), .B0(n7215), .C0(n7214), .Y(n3045)
         );
  AOI2BB2XL U7209 ( .B0(n7303), .B1(n8290), .A0N(n8290), .A1N(image_data[237]), 
        .Y(n7214) );
  AOI22XL U7210 ( .A0(n3357), .A1(n8362), .B0(n8287), .B1(n7078), .Y(n7213) );
  AOI211XL U7211 ( .A0(n3352), .A1(n8293), .B0(n7696), .C0(n7695), .Y(n3046)
         );
  AOI2BB2XL U7212 ( .B0(n3345), .B1(n8290), .A0N(n8290), .A1N(image_data[238]), 
        .Y(n7695) );
  AOI22XL U7213 ( .A0(n8362), .A1(n3353), .B0(n8287), .B1(n3350), .Y(n7694) );
  AOI211XL U7214 ( .A0(n3362), .A1(n8293), .B0(n6716), .C0(n6715), .Y(n3047)
         );
  AOI2BB2XL U7215 ( .B0(n6959), .B1(n8290), .A0N(n8290), .A1N(image_data[239]), 
        .Y(n6715) );
  AOI22XL U7216 ( .A0(n3354), .A1(n8362), .B0(n8287), .B1(n6651), .Y(n6713) );
  AOI211XL U7217 ( .A0(n3355), .A1(n3426), .B0(n7410), .C0(n7409), .Y(n3048)
         );
  AOI2BB2XL U7218 ( .B0(n3367), .B1(n8235), .A0N(n8235), .A1N(image_data[240]), 
        .Y(n7409) );
  AOI22XL U7219 ( .A0(n8114), .A1(n8287), .B0(n8315), .B1(n3360), .Y(n7408) );
  AOI211XL U7220 ( .A0(n3351), .A1(n3426), .B0(n7169), .C0(n7168), .Y(n3049)
         );
  AOI2BB2XL U7221 ( .B0(n3346), .B1(n8235), .A0N(n8235), .A1N(image_data[241]), 
        .Y(n7168) );
  AOI22XL U7222 ( .A0(n7298), .A1(n8287), .B0(n8315), .B1(n3375), .Y(n7167) );
  AOI211XL U7223 ( .A0(n7795), .A1(n3426), .B0(n7841), .C0(n7840), .Y(n3050)
         );
  AOI2BB2XL U7224 ( .B0(n3348), .B1(n8235), .A0N(n8235), .A1N(image_data[242]), 
        .Y(n7840) );
  AOI22XL U7225 ( .A0(n3358), .A1(n8287), .B0(n8315), .B1(n3395), .Y(n7839) );
  AOI211XL U7226 ( .A0(n3387), .A1(n3426), .B0(n8237), .C0(n8236), .Y(n3051)
         );
  AOI2BB2XL U7227 ( .B0(n3347), .B1(n8235), .A0N(n8235), .A1N(image_data[243]), 
        .Y(n8236) );
  AOI22XL U7228 ( .A0(n3389), .A1(n8287), .B0(n8315), .B1(n3349), .Y(n8234) );
  AOI211XL U7229 ( .A0(n8503), .A1(n3426), .B0(n7419), .C0(n7418), .Y(n3052)
         );
  AOI2BB2XL U7230 ( .B0(n6855), .B1(n8235), .A0N(n8235), .A1N(image_data[244]), 
        .Y(n7418) );
  AOI22XL U7231 ( .A0(n3371), .A1(n8287), .B0(n8315), .B1(n6852), .Y(n7417) );
  AOI211XL U7232 ( .A0(n3361), .A1(n3426), .B0(n7151), .C0(n7150), .Y(n3053)
         );
  AOI2BB2XL U7233 ( .B0(n7303), .B1(n8235), .A0N(n8235), .A1N(image_data[245]), 
        .Y(n7150) );
  AOI22XL U7234 ( .A0(n3357), .A1(n8287), .B0(n8315), .B1(n6979), .Y(n7149) );
  AOI211XL U7235 ( .A0(n3352), .A1(n3426), .B0(n7679), .C0(n7678), .Y(n3054)
         );
  AOI2BB2XL U7236 ( .B0(n3345), .B1(n8235), .A0N(n8235), .A1N(image_data[246]), 
        .Y(n7678) );
  AOI22XL U7237 ( .A0(n8287), .A1(n3353), .B0(n8315), .B1(n7581), .Y(n7677) );
  AOI211XL U7238 ( .A0(n3362), .A1(n3426), .B0(n6645), .C0(n6644), .Y(n3055)
         );
  AOI2BB2XL U7239 ( .B0(n6959), .B1(n8235), .A0N(n8235), .A1N(image_data[247]), 
        .Y(n6644) );
  AOI22XL U7240 ( .A0(n3354), .A1(n8287), .B0(n8315), .B1(n6787), .Y(n6642) );
  AOI211XL U7241 ( .A0(n3355), .A1(n8361), .B0(n7532), .C0(n7531), .Y(n3056)
         );
  AOI2BB2XL U7242 ( .B0(n3344), .B1(n8358), .A0N(n8358), .A1N(image_data[248]), 
        .Y(n7531) );
  AOI22XL U7243 ( .A0(n8356), .A1(n3360), .B0(n3378), .B1(n3356), .Y(n7530) );
  AOI211XL U7244 ( .A0(n3351), .A1(n8361), .B0(n7276), .C0(n7275), .Y(n3057)
         );
  AOI2BB2XL U7245 ( .B0(n3346), .B1(n8358), .A0N(n8358), .A1N(image_data[249]), 
        .Y(n7275) );
  AOI22XL U7246 ( .A0(n8356), .A1(n3375), .B0(n3378), .B1(n6332), .Y(n7274) );
  AOI211XL U7247 ( .A0(n7795), .A1(n8361), .B0(n7913), .C0(n7912), .Y(n3058)
         );
  AOI2BB2XL U7248 ( .B0(n3348), .B1(n8358), .A0N(n8358), .A1N(image_data[250]), 
        .Y(n7912) );
  AOI22XL U7249 ( .A0(n3378), .A1(n6880), .B0(n8356), .B1(n3395), .Y(n7911) );
  AOI211XL U7250 ( .A0(n3387), .A1(n8361), .B0(n8360), .C0(n8359), .Y(n3059)
         );
  AOI2BB2XL U7251 ( .B0(n3347), .B1(n8358), .A0N(n8358), .A1N(image_data[251]), 
        .Y(n8359) );
  AOI22XL U7252 ( .A0(n3378), .A1(n6291), .B0(n8356), .B1(n3349), .Y(n8357) );
  AOI211XL U7253 ( .A0(n8503), .A1(n8361), .B0(n7535), .C0(n7534), .Y(n3060)
         );
  AOI2BB2XL U7254 ( .B0(n6855), .B1(n8358), .A0N(n8358), .A1N(image_data[252]), 
        .Y(n7534) );
  AOI22XL U7255 ( .A0(n8356), .A1(n3388), .B0(n3378), .B1(n7326), .Y(n7533) );
  AOI211XL U7256 ( .A0(n3361), .A1(n8361), .B0(n7279), .C0(n7278), .Y(n3061)
         );
  AOI2BB2XL U7257 ( .B0(n7303), .B1(n8358), .A0N(n8358), .A1N(image_data[253]), 
        .Y(n7278) );
  AOI22XL U7258 ( .A0(n8356), .A1(n6979), .B0(n3378), .B1(n7078), .Y(n7277) );
  AOI211XL U7259 ( .A0(n3352), .A1(n8361), .B0(n7735), .C0(n7734), .Y(n3062)
         );
  AOI2BB2XL U7260 ( .B0(n3345), .B1(n8358), .A0N(n8358), .A1N(image_data[254]), 
        .Y(n7734) );
  AOI22XL U7261 ( .A0(n8356), .A1(n7581), .B0(n3378), .B1(n3350), .Y(n7733) );
  AOI211XL U7262 ( .A0(n3362), .A1(n8361), .B0(n6765), .C0(n6764), .Y(n3063)
         );
  AOI2BB2XL U7263 ( .B0(n6959), .B1(n8358), .A0N(n8358), .A1N(image_data[255]), 
        .Y(n6764) );
  AOI22XL U7264 ( .A0(n3378), .A1(n6651), .B0(n8356), .B1(n6787), .Y(n6762) );
  AOI211XL U7265 ( .A0(n3355), .A1(n8258), .B0(n7428), .C0(n7427), .Y(n3064)
         );
  AOI2BB2XL U7266 ( .B0(n3344), .B1(n8255), .A0N(n8255), .A1N(image_data[256]), 
        .Y(n7427) );
  AOI22XL U7267 ( .A0(n8114), .A1(n3378), .B0(n3380), .B1(n3360), .Y(n7426) );
  AOI211XL U7268 ( .A0(n3351), .A1(n8258), .B0(n7181), .C0(n7180), .Y(n3065)
         );
  AOI2BB2XL U7269 ( .B0(n3346), .B1(n8255), .A0N(n8255), .A1N(image_data[257]), 
        .Y(n7180) );
  AOI22XL U7270 ( .A0(n7298), .A1(n3378), .B0(n3380), .B1(n3375), .Y(n7179) );
  AOI211XL U7271 ( .A0(n7795), .A1(n8258), .B0(n7856), .C0(n7855), .Y(n3066)
         );
  AOI2BB2XL U7272 ( .B0(n3348), .B1(n8255), .A0N(n8255), .A1N(image_data[258]), 
        .Y(n7855) );
  AOI22XL U7273 ( .A0(n7923), .A1(n3378), .B0(n3380), .B1(n3395), .Y(n7854) );
  AOI211XL U7274 ( .A0(n3387), .A1(n8258), .B0(n8257), .C0(n8256), .Y(n3067)
         );
  AOI2BB2XL U7275 ( .B0(n3347), .B1(n8255), .A0N(n8255), .A1N(image_data[259]), 
        .Y(n8256) );
  AOI22XL U7276 ( .A0(n3389), .A1(n3378), .B0(n3380), .B1(n3349), .Y(n8254) );
  AOI211XL U7277 ( .A0(n8503), .A1(n8258), .B0(n7425), .C0(n7424), .Y(n3068)
         );
  AOI2BB2XL U7278 ( .B0(n6855), .B1(n8255), .A0N(n8255), .A1N(image_data[260]), 
        .Y(n7424) );
  AOI22XL U7279 ( .A0(n3371), .A1(n3378), .B0(n3380), .B1(n3388), .Y(n7423) );
  AOI21XL U7280 ( .A0(n7898), .A1(n7078), .B0(n6345), .Y(n3069) );
  AOI2BB2XL U7281 ( .B0(n6344), .B1(n8255), .A0N(n8255), .A1N(image_data[261]), 
        .Y(n6345) );
  OAI22XL U7282 ( .A0(n7307), .A1(n6677), .B0(n3391), .B1(n6341), .Y(n6342) );
  AOI211XL U7283 ( .A0(n3352), .A1(n8258), .B0(n7682), .C0(n7681), .Y(n3070)
         );
  AOI2BB2XL U7284 ( .B0(n3345), .B1(n8255), .A0N(n8255), .A1N(image_data[262]), 
        .Y(n7681) );
  AOI22XL U7285 ( .A0(n3378), .A1(n3353), .B0(n3380), .B1(n7581), .Y(n7680) );
  AOI211XL U7286 ( .A0(n3362), .A1(n8258), .B0(n6681), .C0(n6680), .Y(n3071)
         );
  AOI2BB2XL U7287 ( .B0(n6959), .B1(n8255), .A0N(n8255), .A1N(image_data[263]), 
        .Y(n6680) );
  AOI22XL U7288 ( .A0(n3354), .A1(n3378), .B0(n3380), .B1(n3368), .Y(n6679) );
  AOI211XL U7289 ( .A0(n3355), .A1(n8355), .B0(n7526), .C0(n7525), .Y(n3072)
         );
  AOI2BB2XL U7290 ( .B0(n3344), .B1(n8352), .A0N(n8352), .A1N(image_data[264]), 
        .Y(n7525) );
  AOI22XL U7291 ( .A0(n3431), .A1(n3360), .B0(n6143), .B1(n3356), .Y(n7524) );
  AOI211XL U7292 ( .A0(n3351), .A1(n8355), .B0(n7260), .C0(n7259), .Y(n3073)
         );
  AOI2BB2XL U7293 ( .B0(n3346), .B1(n8352), .A0N(n8352), .A1N(image_data[265]), 
        .Y(n7259) );
  AOI22XL U7294 ( .A0(n7898), .A1(n7298), .B0(n6143), .B1(n6332), .Y(n7258) );
  AOI211XL U7295 ( .A0(n7795), .A1(n8355), .B0(n7901), .C0(n7900), .Y(n3074)
         );
  AOI2BB2XL U7296 ( .B0(n3348), .B1(n8352), .A0N(n8352), .A1N(image_data[266]), 
        .Y(n7900) );
  AOI22XL U7297 ( .A0(n7923), .A1(n7898), .B0(n6143), .B1(n6880), .Y(n7899) );
  AOI211XL U7298 ( .A0(n3387), .A1(n8355), .B0(n8354), .C0(n8353), .Y(n3075)
         );
  AOI2BB2XL U7299 ( .B0(n3347), .B1(n8352), .A0N(n8352), .A1N(image_data[267]), 
        .Y(n8353) );
  AOI22XL U7300 ( .A0(n6143), .A1(n6291), .B0(n3431), .B1(n3349), .Y(n8350) );
  AOI211XL U7301 ( .A0(n8503), .A1(n8355), .B0(n7523), .C0(n7522), .Y(n3076)
         );
  AOI2BB2XL U7302 ( .B0(n6855), .B1(n8352), .A0N(n8352), .A1N(image_data[268]), 
        .Y(n7522) );
  AOI22XL U7303 ( .A0(n3371), .A1(n7898), .B0(n3431), .B1(n3388), .Y(n7521) );
  AOI211XL U7304 ( .A0(n3361), .A1(n8355), .B0(n7267), .C0(n7266), .Y(n3077)
         );
  AOI2BB2XL U7305 ( .B0(n7303), .B1(n8352), .A0N(n8352), .A1N(image_data[269]), 
        .Y(n7266) );
  AOI22XL U7306 ( .A0(n3357), .A1(n7898), .B0(n6143), .B1(n7078), .Y(n7265) );
  AOI211XL U7307 ( .A0(n3352), .A1(n8355), .B0(n7729), .C0(n7728), .Y(n3078)
         );
  AOI2BB2XL U7308 ( .B0(n3345), .B1(n8352), .A0N(n8352), .A1N(image_data[270]), 
        .Y(n7728) );
  AOI22XL U7309 ( .A0(n7898), .A1(n3353), .B0(n6143), .B1(n3350), .Y(n7727) );
  AOI211XL U7310 ( .A0(n3362), .A1(n8355), .B0(n6754), .C0(n6753), .Y(n3079)
         );
  AOI2BB2XL U7311 ( .B0(n6959), .B1(n8352), .A0N(n8352), .A1N(image_data[271]), 
        .Y(n6753) );
  AOI22XL U7312 ( .A0(n3354), .A1(n7898), .B0(n6143), .B1(n6651), .Y(n6751) );
  AOI211XL U7313 ( .A0(n3355), .A1(n7929), .B0(n7556), .C0(n7555), .Y(n3080)
         );
  AOI2BB2XL U7314 ( .B0(n3367), .B1(n7926), .A0N(n7926), .A1N(image_data[272]), 
        .Y(n7555) );
  AOI22XL U7315 ( .A0(n8114), .A1(n6143), .B0(n8308), .B1(n3360), .Y(n7554) );
  AOI211XL U7316 ( .A0(n3351), .A1(n7929), .B0(n7301), .C0(n7300), .Y(n3081)
         );
  AOI2BB2XL U7317 ( .B0(n3346), .B1(n7926), .A0N(n7926), .A1N(image_data[273]), 
        .Y(n7300) );
  AOI22XL U7318 ( .A0(n7298), .A1(n6143), .B0(n8308), .B1(n3375), .Y(n7299) );
  AOI211XL U7319 ( .A0(n7795), .A1(n7929), .B0(n7928), .C0(n7927), .Y(n3082)
         );
  AOI2BB2XL U7320 ( .B0(n3348), .B1(n7926), .A0N(n7926), .A1N(image_data[274]), 
        .Y(n7927) );
  AOI22XL U7321 ( .A0(n7923), .A1(n6143), .B0(n8501), .B1(n6880), .Y(n7924) );
  AOI21XL U7322 ( .A0(n8308), .A1(n3349), .B0(n6377), .Y(n3083) );
  AOI2BB2XL U7323 ( .B0(n6376), .B1(n7926), .A0N(n7926), .A1N(image_data[275]), 
        .Y(n6377) );
  AOI211XL U7324 ( .A0(n6143), .A1(n3389), .B0(n6403), .C0(n6373), .Y(n6376)
         );
  AOI211XL U7325 ( .A0(n8503), .A1(n7929), .B0(n7559), .C0(n7558), .Y(n3084)
         );
  AOI2BB2XL U7326 ( .B0(n6855), .B1(n7926), .A0N(n7926), .A1N(image_data[276]), 
        .Y(n7558) );
  AOI22XL U7327 ( .A0(n3371), .A1(n6143), .B0(n8501), .B1(n7326), .Y(n7557) );
  AOI211XL U7328 ( .A0(n3361), .A1(n7929), .B0(n7305), .C0(n7304), .Y(n3085)
         );
  AOI2BB2XL U7329 ( .B0(n7303), .B1(n7926), .A0N(n7926), .A1N(image_data[277]), 
        .Y(n7304) );
  AOI22XL U7330 ( .A0(n3357), .A1(n6143), .B0(n8308), .B1(n6979), .Y(n7302) );
  AOI211XL U7331 ( .A0(n3352), .A1(n7929), .B0(n7745), .C0(n7744), .Y(n3086)
         );
  AOI2BB2XL U7332 ( .B0(n3345), .B1(n7926), .A0N(n7926), .A1N(image_data[278]), 
        .Y(n7744) );
  AOI22XL U7333 ( .A0(n6143), .A1(n3353), .B0(n8308), .B1(n7581), .Y(n7743) );
  AOI211XL U7334 ( .A0(n3362), .A1(n7929), .B0(n6790), .C0(n6789), .Y(n3087)
         );
  AOI2BB2XL U7335 ( .B0(n6959), .B1(n7926), .A0N(n7926), .A1N(image_data[279]), 
        .Y(n6789) );
  AOI22XL U7336 ( .A0(n3354), .A1(n6143), .B0(n8308), .B1(n6787), .Y(n6788) );
  AOI211XL U7337 ( .A0(n3355), .A1(n7910), .B0(n7529), .C0(n7528), .Y(n3088)
         );
  AOI2BB2XL U7338 ( .B0(n3344), .B1(n8507), .A0N(n8507), .A1N(image_data[280]), 
        .Y(n7528) );
  AOI22XL U7339 ( .A0(n8114), .A1(n8501), .B0(n5908), .B1(n3360), .Y(n7527) );
  AOI211XL U7340 ( .A0(n3351), .A1(n7910), .B0(n7273), .C0(n7272), .Y(n3089)
         );
  AOI2BB2XL U7341 ( .B0(n3346), .B1(n8507), .A0N(n8507), .A1N(image_data[281]), 
        .Y(n7272) );
  AOI22XL U7342 ( .A0(n5908), .A1(n3375), .B0(n8499), .B1(n6332), .Y(n7271) );
  AOI211XL U7343 ( .A0(n7795), .A1(n7910), .B0(n7909), .C0(n7908), .Y(n3090)
         );
  AOI2BB2XL U7344 ( .B0(n3348), .B1(n8507), .A0N(n8507), .A1N(image_data[282]), 
        .Y(n7908) );
  AOI22XL U7345 ( .A0(n8499), .A1(n6880), .B0(n5908), .B1(n3395), .Y(n7906) );
  AOI21XL U7346 ( .A0(n3369), .A1(n7910), .B0(n6280), .Y(n3091) );
  AOI22XL U7347 ( .A0(n8499), .A1(n6291), .B0(n5908), .B1(n3349), .Y(n6277) );
  NAND4XL U7348 ( .A(n6855), .B(n8505), .C(n8504), .D(n8507), .Y(n8506) );
  AOI22XL U7349 ( .A0(n5908), .A1(n3388), .B0(n8499), .B1(n7326), .Y(n8505) );
  AOI22XL U7350 ( .A0(n8503), .A1(n8502), .B0(n3371), .B1(n8501), .Y(n8504) );
  AOI211XL U7351 ( .A0(n3361), .A1(n7910), .B0(n7270), .C0(n7269), .Y(n3093)
         );
  AOI2BB2XL U7352 ( .B0(n7303), .B1(n8507), .A0N(n8507), .A1N(image_data[285]), 
        .Y(n7269) );
  AOI22XL U7353 ( .A0(n5908), .A1(n6979), .B0(n8499), .B1(n7078), .Y(n7268) );
  AOI211XL U7354 ( .A0(n3352), .A1(n7910), .B0(n7732), .C0(n7731), .Y(n3094)
         );
  AOI2BB2XL U7355 ( .B0(n3345), .B1(n8507), .A0N(n8507), .A1N(image_data[286]), 
        .Y(n7731) );
  AOI22XL U7356 ( .A0(n8501), .A1(n3353), .B0(n5908), .B1(n7581), .Y(n7730) );
  AOI211XL U7357 ( .A0(n3362), .A1(n7910), .B0(n6757), .C0(n6756), .Y(n3095)
         );
  AOI2BB2XL U7358 ( .B0(n6959), .B1(n8507), .A0N(n8507), .A1N(image_data[287]), 
        .Y(n6756) );
  AOI22XL U7359 ( .A0(n3354), .A1(n8501), .B0(n5908), .B1(n6787), .Y(n6755) );
  AOI211XL U7360 ( .A0(n3355), .A1(n8193), .B0(n7401), .C0(n7400), .Y(n3096)
         );
  AOI2BB2XL U7361 ( .B0(n3344), .B1(n8190), .A0N(n8190), .A1N(image_data[288]), 
        .Y(n7400) );
  AOI22XL U7362 ( .A0(n3381), .A1(n3360), .B0(n7826), .B1(n3356), .Y(n7399) );
  AOI211XL U7363 ( .A0(n3351), .A1(n8193), .B0(n7142), .C0(n7141), .Y(n3097)
         );
  AOI2BB2XL U7364 ( .B0(n3346), .B1(n8190), .A0N(n8190), .A1N(image_data[289]), 
        .Y(n7141) );
  AOI22XL U7365 ( .A0(n7298), .A1(n8499), .B0(n3381), .B1(n3375), .Y(n7140) );
  AOI211XL U7366 ( .A0(n7795), .A1(n8193), .B0(n7829), .C0(n7828), .Y(n3098)
         );
  AOI2BB2XL U7367 ( .B0(n3348), .B1(n8190), .A0N(n8190), .A1N(image_data[290]), 
        .Y(n7828) );
  AOI22XL U7368 ( .A0(n7826), .A1(n6880), .B0(n3381), .B1(n3395), .Y(n7827) );
  AOI211XL U7369 ( .A0(n3387), .A1(n8193), .B0(n8192), .C0(n8191), .Y(n3099)
         );
  AOI2BB2XL U7370 ( .B0(n3347), .B1(n8190), .A0N(n8190), .A1N(image_data[291]), 
        .Y(n8191) );
  AOI22XL U7371 ( .A0(n3389), .A1(n8499), .B0(n3381), .B1(n3349), .Y(n8189) );
  AOI211XL U7372 ( .A0(n8503), .A1(n8193), .B0(n7395), .C0(n7394), .Y(n3100)
         );
  AOI2BB2XL U7373 ( .B0(n6855), .B1(n8190), .A0N(n8190), .A1N(image_data[292]), 
        .Y(n7394) );
  AOI22XL U7374 ( .A0(n3381), .A1(n3388), .B0(n7826), .B1(n7326), .Y(n7393) );
  AOI211XL U7375 ( .A0(n3361), .A1(n8193), .B0(n7157), .C0(n7156), .Y(n3101)
         );
  AOI2BB2XL U7376 ( .B0(n7303), .B1(n8190), .A0N(n8190), .A1N(image_data[293]), 
        .Y(n7156) );
  AOI22XL U7377 ( .A0(n3381), .A1(n6979), .B0(n7826), .B1(n7078), .Y(n7155) );
  AOI211XL U7378 ( .A0(n3352), .A1(n8193), .B0(n7661), .C0(n7660), .Y(n3102)
         );
  AOI2BB2XL U7379 ( .B0(n3345), .B1(n8190), .A0N(n8190), .A1N(image_data[294]), 
        .Y(n7660) );
  AOI22XL U7380 ( .A0(n3381), .A1(n7581), .B0(n7826), .B1(n3350), .Y(n7659) );
  AOI211XL U7381 ( .A0(n3362), .A1(n8193), .B0(n6637), .C0(n6636), .Y(n3103)
         );
  AOI2BB2XL U7382 ( .B0(n6959), .B1(n8190), .A0N(n8190), .A1N(image_data[295]), 
        .Y(n6636) );
  AOI22XL U7383 ( .A0(n3354), .A1(n8499), .B0(n3381), .B1(n3368), .Y(n6635) );
  AOI211XL U7384 ( .A0(n3355), .A1(n7486), .B0(n7485), .C0(n7484), .Y(n3104)
         );
  AOI2BB2XL U7385 ( .B0(n3367), .B1(n7483), .A0N(n7483), .A1N(image_data[296]), 
        .Y(n7484) );
  AOI22XL U7386 ( .A0(n7888), .A1(n3360), .B0(n8315), .B1(n3356), .Y(n7482) );
  AOI211XL U7387 ( .A0(n3351), .A1(n7486), .B0(n7239), .C0(n7238), .Y(n3105)
         );
  AOI2BB2XL U7388 ( .B0(n3346), .B1(n7483), .A0N(n7483), .A1N(image_data[297]), 
        .Y(n7238) );
  AOI22XL U7389 ( .A0(n7888), .A1(n3375), .B0(n8315), .B1(n6332), .Y(n7237) );
  OAI22XL U7390 ( .A0(n7895), .A1(n7878), .B0(n7773), .B1(n8289), .Y(n6397) );
  AOI2BB2XL U7391 ( .B0(n6395), .B1(n7483), .A0N(n7483), .A1N(image_data[298]), 
        .Y(n6396) );
  AOI221XL U7392 ( .A0(image_data[299]), .A1(n3423), .B0(n6413), .B1(n7483), 
        .C0(n6412), .Y(n3107) );
  AOI22XL U7393 ( .A0(n8315), .A1(n6291), .B0(n7888), .B1(n3349), .Y(n6411) );
  OAI22XL U7394 ( .A0(n3370), .A1(n8136), .B0(n8035), .B1(n8289), .Y(n6394) );
  AOI2BB2XL U7395 ( .B0(n6392), .B1(n7483), .A0N(n7483), .A1N(image_data[300]), 
        .Y(n6393) );
  AOI211XL U7396 ( .A0(n3361), .A1(n7486), .B0(n7242), .C0(n7241), .Y(n3109)
         );
  AOI2BB2XL U7397 ( .B0(n7303), .B1(n7483), .A0N(n7483), .A1N(image_data[301]), 
        .Y(n7241) );
  AOI22XL U7398 ( .A0(n7888), .A1(n6979), .B0(n8315), .B1(n7078), .Y(n7240) );
  AOI221XL U7399 ( .A0(image_data[302]), .A1(n3423), .B0(n6954), .B1(n7483), 
        .C0(n6953), .Y(n3110) );
  AOI22XL U7400 ( .A0(n7888), .A1(n7581), .B0(n8315), .B1(n3350), .Y(n6952) );
  AOI211XL U7401 ( .A0(n3423), .A1(image_data[303]), .B0(n6967), .C0(n6966), 
        .Y(n3111) );
  OAI22XL U7402 ( .A0(n7570), .A1(n7878), .B0(n3394), .B1(n8136), .Y(n6966) );
  AOI21XL U7403 ( .A0(n6959), .A1(n6965), .B0(n3423), .Y(n6967) );
  AOI22XL U7404 ( .A0(n3362), .A1(n6964), .B0(n6973), .B1(n7826), .Y(n6965) );
  AOI211XL U7405 ( .A0(n3355), .A1(n8321), .B0(n7496), .C0(n7495), .Y(n3112)
         );
  AOI2BB2XL U7406 ( .B0(n3344), .B1(n8318), .A0N(n8318), .A1N(image_data[304]), 
        .Y(n7495) );
  AOI22XL U7407 ( .A0(n8315), .A1(n8114), .B0(n8356), .B1(n3356), .Y(n7494) );
  AOI211XL U7408 ( .A0(n3351), .A1(n8321), .B0(n7254), .C0(n7253), .Y(n3113)
         );
  AOI2BB2XL U7409 ( .B0(n3366), .B1(n8318), .A0N(n8318), .A1N(image_data[305]), 
        .Y(n7253) );
  AOI22XL U7410 ( .A0(n8315), .A1(n7298), .B0(n8356), .B1(n6332), .Y(n7252) );
  AOI211XL U7411 ( .A0(n7795), .A1(n8321), .B0(n7880), .C0(n7879), .Y(n3114)
         );
  AOI2BB2XL U7412 ( .B0(n3348), .B1(n8318), .A0N(n8318), .A1N(image_data[306]), 
        .Y(n7879) );
  AOI22XL U7413 ( .A0(n8356), .A1(n6880), .B0(n7887), .B1(n3395), .Y(n7877) );
  AOI211XL U7414 ( .A0(n3387), .A1(n8321), .B0(n8320), .C0(n8319), .Y(n3115)
         );
  AOI2BB2XL U7415 ( .B0(n3347), .B1(n8318), .A0N(n8318), .A1N(image_data[307]), 
        .Y(n8319) );
  AOI22XL U7416 ( .A0(n3389), .A1(n8315), .B0(n8356), .B1(n6291), .Y(n8316) );
  AOI211XL U7417 ( .A0(n8321), .A1(n8503), .B0(n7061), .C0(n7060), .Y(n3116)
         );
  NOR2XL U7418 ( .A(n3370), .B(n8317), .Y(n7061) );
  AOI32XL U7419 ( .A0(n6855), .A1(n8318), .A2(n7059), .B0(n3412), .B1(n8536), 
        .Y(n7060) );
  AOI22XL U7420 ( .A0(n3371), .A1(n8315), .B0(n8356), .B1(n7326), .Y(n7059) );
  AOI211XL U7421 ( .A0(n3361), .A1(n8321), .B0(n7251), .C0(n7250), .Y(n3117)
         );
  AOI2BB2XL U7422 ( .B0(n7303), .B1(n8318), .A0N(n8318), .A1N(image_data[309]), 
        .Y(n7250) );
  AOI22XL U7423 ( .A0(n7938), .A1(n8315), .B0(n7887), .B1(n6979), .Y(n7249) );
  AOI211XL U7424 ( .A0(n3352), .A1(n8321), .B0(n7716), .C0(n7715), .Y(n3118)
         );
  AOI2BB2XL U7425 ( .B0(n3345), .B1(n8318), .A0N(n8318), .A1N(image_data[310]), 
        .Y(n7715) );
  AOI22XL U7426 ( .A0(n8315), .A1(n3353), .B0(n7887), .B1(n7581), .Y(n7714) );
  AOI211XL U7427 ( .A0(n3362), .A1(n8321), .B0(n6732), .C0(n6731), .Y(n3119)
         );
  AOI2BB2XL U7428 ( .B0(n6959), .B1(n8318), .A0N(n8318), .A1N(image_data[311]), 
        .Y(n6731) );
  AOI22XL U7429 ( .A0(n3354), .A1(n8315), .B0(n7887), .B1(n3368), .Y(n6730) );
  AOI221XL U7430 ( .A0(image_data[312]), .A1(n8026), .B0(n6997), .B1(n8131), 
        .C0(n6996), .Y(n3120) );
  AOI22XL U7431 ( .A0(n8356), .A1(n8114), .B0(n3380), .B1(n3356), .Y(n6995) );
  AOI211XL U7432 ( .A0(n3351), .A1(n8134), .B0(n7064), .C0(n7063), .Y(n3121)
         );
  AOI2BB2XL U7433 ( .B0(n3366), .B1(n8131), .A0N(n8131), .A1N(image_data[313]), 
        .Y(n7063) );
  AOI22XL U7434 ( .A0(n3455), .A1(n3375), .B0(n3380), .B1(n6332), .Y(n7062) );
  AOI211XL U7435 ( .A0(n7795), .A1(n8134), .B0(n7794), .C0(n7793), .Y(n3122)
         );
  AOI2BB2XL U7436 ( .B0(n3348), .B1(n8131), .A0N(n8131), .A1N(image_data[314]), 
        .Y(n7793) );
  AOI22XL U7437 ( .A0(n3380), .A1(n6880), .B0(n3455), .B1(n3395), .Y(n7792) );
  AOI211XL U7438 ( .A0(n3387), .A1(n8134), .B0(n8133), .C0(n8132), .Y(n3123)
         );
  AOI2BB2XL U7439 ( .B0(n3347), .B1(n8131), .A0N(n8131), .A1N(image_data[315]), 
        .Y(n8132) );
  AOI22XL U7440 ( .A0(n3380), .A1(n6291), .B0(n3455), .B1(n3349), .Y(n8129) );
  AOI211XL U7441 ( .A0(n8026), .A1(image_data[316]), .B0(n8025), .C0(n8024), 
        .Y(n3124) );
  OAI22XL U7442 ( .A0(n3370), .A1(n8023), .B0(n8035), .B1(n8130), .Y(n8024) );
  AOI21XL U7443 ( .A0(n6855), .A1(n8022), .B0(n8026), .Y(n8025) );
  AOI22XL U7444 ( .A0(n8503), .A1(n8021), .B0(n3380), .B1(n7326), .Y(n8022) );
  AOI211XL U7445 ( .A0(n3361), .A1(n8134), .B0(n7067), .C0(n7066), .Y(n3125)
         );
  AOI2BB2XL U7446 ( .B0(n7303), .B1(n8131), .A0N(n8131), .A1N(image_data[317]), 
        .Y(n7066) );
  AOI22XL U7447 ( .A0(n3455), .A1(n6979), .B0(n3380), .B1(n7078), .Y(n7065) );
  AOI211XL U7448 ( .A0(n3352), .A1(n8134), .B0(n7628), .C0(n7627), .Y(n3126)
         );
  AOI2BB2XL U7449 ( .B0(n3345), .B1(n8131), .A0N(n8131), .A1N(image_data[318]), 
        .Y(n7627) );
  AOI22XL U7450 ( .A0(n3455), .A1(n7581), .B0(n3380), .B1(n3350), .Y(n7626) );
  AOI221XL U7451 ( .A0(image_data[319]), .A1(n8026), .B0(n7580), .B1(n8131), 
        .C0(n7579), .Y(n3127) );
  AOI22XL U7452 ( .A0(n3380), .A1(n6651), .B0(n3455), .B1(n3368), .Y(n7576) );
  AOI211XL U7453 ( .A0(n3355), .A1(n8169), .B0(n7358), .C0(n7357), .Y(n3128)
         );
  AOI2BB2XL U7454 ( .B0(n3344), .B1(n8166), .A0N(n8166), .A1N(image_data[320]), 
        .Y(n7357) );
  AOI22XL U7455 ( .A0(n3380), .A1(n8114), .B0(n3431), .B1(n3356), .Y(n7356) );
  AOI211XL U7456 ( .A0(n3351), .A1(n8169), .B0(n7093), .C0(n7092), .Y(n3129)
         );
  AOI2BB2XL U7457 ( .B0(n3366), .B1(n8166), .A0N(n8166), .A1N(image_data[321]), 
        .Y(n7092) );
  AOI22XL U7458 ( .A0(n3380), .A1(n7298), .B0(n3431), .B1(n6332), .Y(n7091) );
  AOI211XL U7459 ( .A0(n7795), .A1(n8169), .B0(n7819), .C0(n7818), .Y(n3130)
         );
  AOI2BB2XL U7460 ( .B0(n3348), .B1(n8166), .A0N(n8166), .A1N(image_data[322]), 
        .Y(n7818) );
  AOI22XL U7461 ( .A0(n7923), .A1(n3380), .B0(n3431), .B1(n6880), .Y(n7817) );
  AOI211XL U7462 ( .A0(n3387), .A1(n8169), .B0(n8168), .C0(n8167), .Y(n3131)
         );
  AOI2BB2XL U7463 ( .B0(n3347), .B1(n8166), .A0N(n8166), .A1N(image_data[323]), 
        .Y(n8167) );
  AOI22XL U7464 ( .A0(n3389), .A1(n3380), .B0(n3431), .B1(n6291), .Y(n8164) );
  AOI211XL U7465 ( .A0(n8503), .A1(n8169), .B0(n7341), .C0(n7340), .Y(n3132)
         );
  AOI2BB2XL U7466 ( .B0(n6855), .B1(n8166), .A0N(n8166), .A1N(image_data[324]), 
        .Y(n7340) );
  AOI22XL U7467 ( .A0(n3371), .A1(n3380), .B0(n3431), .B1(n7326), .Y(n7339) );
  AOI211XL U7468 ( .A0(n3361), .A1(n8169), .B0(n7090), .C0(n7089), .Y(n3133)
         );
  AOI2BB2XL U7469 ( .B0(n7303), .B1(n8166), .A0N(n8166), .A1N(image_data[325]), 
        .Y(n7089) );
  AOI22XL U7470 ( .A0(n7938), .A1(n3380), .B0(n3431), .B1(n7078), .Y(n7088) );
  AOI21XL U7471 ( .A0(n3352), .A1(n8169), .B0(n6171), .Y(n3134) );
  AOI22XL U7472 ( .A0(n8238), .A1(n7581), .B0(n3431), .B1(n3350), .Y(n6168) );
  AOI211XL U7473 ( .A0(n3362), .A1(n8169), .B0(n6601), .C0(n6600), .Y(n3135)
         );
  AOI2BB2XL U7474 ( .B0(n6959), .B1(n8166), .A0N(n8166), .A1N(image_data[327]), 
        .Y(n6600) );
  AOI22XL U7475 ( .A0(n3354), .A1(n3380), .B0(n3431), .B1(n6651), .Y(n6599) );
  AOI211XL U7476 ( .A0(n3355), .A1(n8314), .B0(n7499), .C0(n7498), .Y(n3136)
         );
  AOI2BB2XL U7477 ( .B0(n3344), .B1(n8311), .A0N(n8311), .A1N(image_data[328]), 
        .Y(n7498) );
  AOI22XL U7478 ( .A0(n3431), .A1(n8114), .B0(n8308), .B1(n3356), .Y(n7497) );
  AOI211XL U7479 ( .A0(n3351), .A1(n8314), .B0(n7248), .C0(n7247), .Y(n3137)
         );
  AOI2BB2XL U7480 ( .B0(n3366), .B1(n8311), .A0N(n8311), .A1N(image_data[329]), 
        .Y(n7247) );
  AOI22XL U7481 ( .A0(n3431), .A1(n7298), .B0(n8308), .B1(n6943), .Y(n7246) );
  AOI211XL U7482 ( .A0(n7795), .A1(n8314), .B0(n7883), .C0(n7882), .Y(n3138)
         );
  AOI2BB2XL U7483 ( .B0(n3348), .B1(n8311), .A0N(n8311), .A1N(image_data[330]), 
        .Y(n7882) );
  AOI22XL U7484 ( .A0(n7923), .A1(n3431), .B0(n8308), .B1(n6880), .Y(n7881) );
  AOI211XL U7485 ( .A0(n3387), .A1(n8314), .B0(n8313), .C0(n8312), .Y(n3139)
         );
  AOI2BB2XL U7486 ( .B0(n3347), .B1(n8311), .A0N(n8311), .A1N(image_data[331]), 
        .Y(n8312) );
  AOI22XL U7487 ( .A0(n3389), .A1(n3431), .B0(n8308), .B1(n6291), .Y(n8309) );
  AOI211XL U7488 ( .A0(n8503), .A1(n8314), .B0(n7502), .C0(n7501), .Y(n3140)
         );
  AOI2BB2XL U7489 ( .B0(n6855), .B1(n8311), .A0N(n8311), .A1N(image_data[332]), 
        .Y(n7501) );
  AOI22XL U7490 ( .A0(n3371), .A1(n3431), .B0(n8308), .B1(n7326), .Y(n7500) );
  AOI211XL U7491 ( .A0(n8314), .A1(n3361), .B0(n7942), .C0(n7941), .Y(n3141)
         );
  OAI2BB2XL U7492 ( .B0(n7963), .B1(n8310), .A0N(image_data[333]), .A1N(n7940), 
        .Y(n7941) );
  AOI21XL U7493 ( .A0(n8496), .A1(n7939), .B0(n7940), .Y(n7942) );
  AOI22XL U7494 ( .A0(n7938), .A1(n3431), .B0(n8308), .B1(n7078), .Y(n7939) );
  AOI211XL U7495 ( .A0(n3352), .A1(n8314), .B0(n7710), .C0(n7709), .Y(n3142)
         );
  AOI2BB2XL U7496 ( .B0(n3345), .B1(n8311), .A0N(n8311), .A1N(image_data[334]), 
        .Y(n7709) );
  AOI22XL U7497 ( .A0(n3431), .A1(n3353), .B0(n8308), .B1(n3350), .Y(n7708) );
  AOI211XL U7498 ( .A0(n3362), .A1(n8314), .B0(n6738), .C0(n6737), .Y(n3143)
         );
  AOI2BB2XL U7499 ( .B0(n6586), .B1(n8311), .A0N(n8311), .A1N(image_data[335]), 
        .Y(n6737) );
  AOI22XL U7500 ( .A0(n3354), .A1(n3431), .B0(n8308), .B1(n6651), .Y(n6736) );
  AOI21XL U7501 ( .A0(n3373), .A1(n3434), .B0(n6130), .Y(n3144) );
  AOI22XL U7502 ( .A0(n8114), .A1(n8308), .B0(n8214), .B1(n3360), .Y(n6128) );
  AOI211XL U7503 ( .A0(n3351), .A1(n3434), .B0(n7200), .C0(n7199), .Y(n3145)
         );
  AOI2BB2XL U7504 ( .B0(n3366), .B1(n8269), .A0N(n8269), .A1N(image_data[337]), 
        .Y(n7199) );
  AOI22XL U7505 ( .A0(n8308), .A1(n7298), .B0(n5908), .B1(n6332), .Y(n7198) );
  AOI221XL U7506 ( .A0(image_data[338]), .A1(n6884), .B0(n6883), .B1(n8269), 
        .C0(n6882), .Y(n3146) );
  OAI2BB1XL U7507 ( .A0N(n6879), .A1N(n6878), .B0(n3348), .Y(n6883) );
  AOI22XL U7508 ( .A0(n5908), .A1(n6880), .B0(n8214), .B1(n3395), .Y(n6881) );
  AOI211XL U7509 ( .A0(n3387), .A1(n3434), .B0(n8271), .C0(n8270), .Y(n3147)
         );
  AOI2BB2XL U7510 ( .B0(n3347), .B1(n8269), .A0N(n8269), .A1N(image_data[339]), 
        .Y(n8270) );
  AOI22XL U7511 ( .A0(n3389), .A1(n8308), .B0(n5908), .B1(n6291), .Y(n8266) );
  AOI211XL U7512 ( .A0(n8503), .A1(n3434), .B0(n7453), .C0(n7452), .Y(n3148)
         );
  AOI2BB2XL U7513 ( .B0(n6855), .B1(n8269), .A0N(n8269), .A1N(image_data[340]), 
        .Y(n7452) );
  AOI22XL U7514 ( .A0(n3371), .A1(n8308), .B0(n5908), .B1(n7326), .Y(n7451) );
  AOI211XL U7515 ( .A0(n3361), .A1(n3434), .B0(n7197), .C0(n7196), .Y(n3149)
         );
  AOI2BB2XL U7516 ( .B0(n7303), .B1(n8269), .A0N(n8269), .A1N(image_data[341]), 
        .Y(n7196) );
  AOI22XL U7517 ( .A0(n3357), .A1(n8308), .B0(n5908), .B1(n7078), .Y(n7195) );
  AOI21XL U7518 ( .A0(n3352), .A1(n3434), .B0(n6158), .Y(n3150) );
  AOI22XL U7519 ( .A0(n8308), .A1(n3353), .B0(n5908), .B1(n3350), .Y(n6156) );
  AOI211XL U7520 ( .A0(n3362), .A1(n3434), .B0(n6696), .C0(n6695), .Y(n3151)
         );
  AOI2BB2XL U7521 ( .B0(n6959), .B1(n8269), .A0N(n8269), .A1N(image_data[343]), 
        .Y(n6695) );
  AOI22XL U7522 ( .A0(n3354), .A1(n8308), .B0(n5908), .B1(n6651), .Y(n6694) );
  AOI211XL U7523 ( .A0(n3373), .A1(n8163), .B0(n7361), .C0(n7360), .Y(n3152)
         );
  AOI2BB2XL U7524 ( .B0(n3344), .B1(n8160), .A0N(n8160), .A1N(image_data[344]), 
        .Y(n7360) );
  AOI22XL U7525 ( .A0(n5908), .A1(n8114), .B0(n3381), .B1(n3356), .Y(n7359) );
  AOI211XL U7526 ( .A0(n3351), .A1(n8163), .B0(n7109), .C0(n7108), .Y(n3153)
         );
  AOI2BB2XL U7527 ( .B0(n3366), .B1(n8160), .A0N(n8160), .A1N(image_data[345]), 
        .Y(n7108) );
  AOI22XL U7528 ( .A0(n5908), .A1(n7298), .B0(n3381), .B1(n6332), .Y(n7107) );
  AOI21XL U7529 ( .A0(n7795), .A1(n8163), .B0(n5913), .Y(n3154) );
  AOI22XL U7530 ( .A0(n7923), .A1(n5908), .B0(n3381), .B1(n6880), .Y(n5911) );
  AOI211XL U7531 ( .A0(n3387), .A1(n8163), .B0(n8162), .C0(n8161), .Y(n3155)
         );
  AOI2BB2XL U7532 ( .B0(n3347), .B1(n8160), .A0N(n8160), .A1N(image_data[347]), 
        .Y(n8161) );
  AOI22XL U7533 ( .A0(n3389), .A1(n5908), .B0(n3381), .B1(n6291), .Y(n8158) );
  AOI211XL U7534 ( .A0(n8503), .A1(n8163), .B0(n7355), .C0(n7354), .Y(n3156)
         );
  AOI2BB2XL U7535 ( .B0(n6855), .B1(n8160), .A0N(n8160), .A1N(image_data[348]), 
        .Y(n7354) );
  AOI22XL U7536 ( .A0(n3371), .A1(n5908), .B0(n3381), .B1(n7326), .Y(n7353) );
  AOI211XL U7537 ( .A0(n8163), .A1(n3361), .B0(n7937), .C0(n7936), .Y(n3157)
         );
  OAI2BB2XL U7538 ( .B0(n7963), .B1(n8159), .A0N(image_data[349]), .A1N(n7935), 
        .Y(n7936) );
  AOI21XL U7539 ( .A0(n8496), .A1(n7934), .B0(n7935), .Y(n7937) );
  AOI22XL U7540 ( .A0(n3357), .A1(n5908), .B0(n3381), .B1(n7078), .Y(n7934) );
  AOI211XL U7541 ( .A0(n3352), .A1(n8163), .B0(n7646), .C0(n7645), .Y(n3158)
         );
  AOI2BB2XL U7542 ( .B0(n3345), .B1(n8160), .A0N(n8160), .A1N(image_data[350]), 
        .Y(n7645) );
  AOI22XL U7543 ( .A0(n5908), .A1(n3353), .B0(n3381), .B1(n3350), .Y(n7644) );
  AOI211XL U7544 ( .A0(n3362), .A1(n8163), .B0(n6610), .C0(n6609), .Y(n3159)
         );
  AOI2BB2XL U7545 ( .B0(n6959), .B1(n8160), .A0N(n8160), .A1N(image_data[351]), 
        .Y(n6609) );
  AOI22XL U7546 ( .A0(n3354), .A1(n5908), .B0(n3381), .B1(n6651), .Y(n6608) );
  AOI211XL U7547 ( .A0(n3373), .A1(n8140), .B0(n7322), .C0(n7321), .Y(n3160)
         );
  AOI2BB2XL U7548 ( .B0(n3344), .B1(n8137), .A0N(n8137), .A1N(image_data[352]), 
        .Y(n7321) );
  AOI22XL U7549 ( .A0(n8114), .A1(n3381), .B0(n3452), .B1(n3360), .Y(n7320) );
  AOI211XL U7550 ( .A0(n3351), .A1(n8140), .B0(n7071), .C0(n7070), .Y(n3161)
         );
  AOI2BB2XL U7551 ( .B0(n3366), .B1(n8137), .A0N(n8137), .A1N(image_data[353]), 
        .Y(n7070) );
  AOI22XL U7552 ( .A0(n7298), .A1(n3381), .B0(n3452), .B1(n3375), .Y(n7069) );
  AOI211XL U7553 ( .A0(n7795), .A1(n8140), .B0(n7804), .C0(n7803), .Y(n3162)
         );
  AOI2BB2XL U7554 ( .B0(n3348), .B1(n8137), .A0N(n8137), .A1N(image_data[354]), 
        .Y(n7803) );
  AOI22XL U7555 ( .A0(n7923), .A1(n3381), .B0(n3452), .B1(n3395), .Y(n7802) );
  AOI211XL U7556 ( .A0(n3387), .A1(n8140), .B0(n8139), .C0(n8138), .Y(n3163)
         );
  AOI2BB2XL U7557 ( .B0(n3347), .B1(n8137), .A0N(n8137), .A1N(image_data[355]), 
        .Y(n8138) );
  AOI22XL U7558 ( .A0(n3389), .A1(n3381), .B0(n3452), .B1(n3349), .Y(n8135) );
  AOI211XL U7559 ( .A0(n8503), .A1(n8140), .B0(n7325), .C0(n7324), .Y(n3164)
         );
  AOI2BB2XL U7560 ( .B0(n6855), .B1(n8137), .A0N(n8137), .A1N(image_data[356]), 
        .Y(n7324) );
  AOI22XL U7561 ( .A0(n3371), .A1(n3381), .B0(n3452), .B1(n3388), .Y(n7323) );
  AOI21XL U7562 ( .A0(n3452), .A1(n6979), .B0(n6328), .Y(n3165) );
  AOI32XL U7563 ( .A0(n6327), .A1(n8137), .A2(n6326), .B0(n6325), .B1(n8535), 
        .Y(n6328) );
  AOI22XL U7564 ( .A0(n7938), .A1(n3381), .B0(n7888), .B1(n7078), .Y(n6327) );
  AOI211XL U7565 ( .A0(n3352), .A1(n8140), .B0(n7640), .C0(n7639), .Y(n3166)
         );
  AOI2BB2XL U7566 ( .B0(n3345), .B1(n8137), .A0N(n8137), .A1N(image_data[358]), 
        .Y(n7639) );
  AOI22XL U7567 ( .A0(n3381), .A1(n3353), .B0(n3452), .B1(n7581), .Y(n7638) );
  AOI211XL U7568 ( .A0(n3362), .A1(n8140), .B0(n6595), .C0(n6594), .Y(n3167)
         );
  AOI2BB2XL U7569 ( .B0(n6959), .B1(n8137), .A0N(n8137), .A1N(image_data[359]), 
        .Y(n6594) );
  AOI22XL U7570 ( .A0(n3354), .A1(n3381), .B0(n3452), .B1(n3368), .Y(n6593) );
  AOI211XL U7571 ( .A0(n3373), .A1(n7893), .B0(n7509), .C0(n7508), .Y(n3168)
         );
  AOI2BB2XL U7572 ( .B0(n3344), .B1(n7890), .A0N(n7890), .A1N(image_data[360]), 
        .Y(n7508) );
  AOI22XL U7573 ( .A0(n7888), .A1(n8114), .B0(n7887), .B1(n3356), .Y(n7506) );
  AOI21XL U7574 ( .A0(n3351), .A1(n7893), .B0(n5703), .Y(n3169) );
  AOI22XL U7575 ( .A0(n7888), .A1(n7298), .B0(n7887), .B1(n6332), .Y(n5701) );
  AOI211XL U7576 ( .A0(n7795), .A1(n7893), .B0(n7892), .C0(n7891), .Y(n3170)
         );
  AOI2BB2XL U7577 ( .B0(n3348), .B1(n7890), .A0N(n7890), .A1N(image_data[362]), 
        .Y(n7891) );
  AOI22XL U7578 ( .A0(n7923), .A1(n7888), .B0(n7887), .B1(n6880), .Y(n7889) );
  AOI21XL U7579 ( .A0(n3369), .A1(n7893), .B0(n6274), .Y(n3171) );
  AOI22XL U7580 ( .A0(n7887), .A1(n6291), .B0(n8492), .B1(n3349), .Y(n6271) );
  AOI211XL U7581 ( .A0(n8503), .A1(n7893), .B0(n7505), .C0(n7504), .Y(n3172)
         );
  AOI2BB2XL U7582 ( .B0(n6855), .B1(n7890), .A0N(n7890), .A1N(image_data[364]), 
        .Y(n7504) );
  AOI22XL U7583 ( .A0(n3371), .A1(n7888), .B0(n7887), .B1(n7326), .Y(n7503) );
  AOI211XL U7584 ( .A0(n3361), .A1(n7893), .B0(n7257), .C0(n7256), .Y(n3173)
         );
  AOI2BB2XL U7585 ( .B0(n8496), .B1(n7890), .A0N(n7890), .A1N(image_data[365]), 
        .Y(n7256) );
  AOI22XL U7586 ( .A0(n8492), .A1(n6979), .B0(n7887), .B1(n7078), .Y(n7255) );
  AOI211XL U7587 ( .A0(n3352), .A1(n7893), .B0(n7719), .C0(n7718), .Y(n3174)
         );
  AOI2BB2XL U7588 ( .B0(n3345), .B1(n7890), .A0N(n7890), .A1N(image_data[366]), 
        .Y(n7718) );
  AOI22XL U7589 ( .A0(n7888), .A1(n3353), .B0(n7887), .B1(n3350), .Y(n7717) );
  AOI211XL U7590 ( .A0(n3362), .A1(n7893), .B0(n6741), .C0(n6740), .Y(n3175)
         );
  AOI2BB2XL U7591 ( .B0(n6959), .B1(n7890), .A0N(n7890), .A1N(image_data[367]), 
        .Y(n6740) );
  AOI22XL U7592 ( .A0(n3354), .A1(n7888), .B0(n7887), .B1(n6651), .Y(n6739) );
  AOI211XL U7593 ( .A0(n3373), .A1(n7701), .B0(n7472), .C0(n7471), .Y(n3176)
         );
  AOI2BB2XL U7594 ( .B0(n3367), .B1(n7698), .A0N(n7698), .A1N(image_data[368]), 
        .Y(n7471) );
  AOI22XL U7595 ( .A0(n7887), .A1(n8114), .B0(n3455), .B1(n3356), .Y(n7470) );
  AOI211XL U7596 ( .A0(n3351), .A1(n7701), .B0(n7224), .C0(n7223), .Y(n3177)
         );
  AOI2BB2XL U7597 ( .B0(n3366), .B1(n7698), .A0N(n7698), .A1N(image_data[369]), 
        .Y(n7223) );
  AOI22XL U7598 ( .A0(n7887), .A1(n7298), .B0(n3455), .B1(n6332), .Y(n7222) );
  AOI21XL U7599 ( .A0(n7795), .A1(n7701), .B0(n5920), .Y(n3178) );
  AOI22XL U7600 ( .A0(n7923), .A1(n7887), .B0(n8490), .B1(n3395), .Y(n5917) );
  AOI21XL U7601 ( .A0(n3369), .A1(n7701), .B0(n6298), .Y(n3179) );
  AOI2BB2XL U7602 ( .B0(n6297), .B1(n7698), .A0N(n7698), .A1N(image_data[371]), 
        .Y(n6298) );
  AOI211XL U7603 ( .A0(n7887), .A1(n3389), .B0(n6403), .C0(n6296), .Y(n6297)
         );
  OAI22XL U7604 ( .A0(n8447), .A1(n8023), .B0(n3386), .B1(n8125), .Y(n6296) );
  AOI211XL U7605 ( .A0(n8503), .A1(n7701), .B0(n7475), .C0(n7474), .Y(n3180)
         );
  AOI2BB2XL U7606 ( .B0(n6855), .B1(n7698), .A0N(n7698), .A1N(image_data[372]), 
        .Y(n7474) );
  AOI22XL U7607 ( .A0(n3371), .A1(n7887), .B0(n3455), .B1(n7326), .Y(n7473) );
  AOI211XL U7608 ( .A0(n3361), .A1(n7701), .B0(n7227), .C0(n7226), .Y(n3181)
         );
  AOI2BB2XL U7609 ( .B0(n7303), .B1(n7698), .A0N(n7698), .A1N(image_data[373]), 
        .Y(n7226) );
  AOI22XL U7610 ( .A0(n3357), .A1(n7887), .B0(n3455), .B1(n7078), .Y(n7225) );
  AOI211XL U7611 ( .A0(n3352), .A1(n7701), .B0(n7700), .C0(n7699), .Y(n3182)
         );
  AOI2BB2XL U7612 ( .B0(n3345), .B1(n7698), .A0N(n7698), .A1N(image_data[374]), 
        .Y(n7699) );
  AOI22XL U7613 ( .A0(n7887), .A1(n3353), .B0(n3455), .B1(n3350), .Y(n7697) );
  AOI211XL U7614 ( .A0(n3362), .A1(n7701), .B0(n6719), .C0(n6718), .Y(n3183)
         );
  AOI2BB2XL U7615 ( .B0(n6959), .B1(n7698), .A0N(n7698), .A1N(image_data[375]), 
        .Y(n6718) );
  AOI22XL U7616 ( .A0(n3354), .A1(n7887), .B0(n3455), .B1(n6651), .Y(n6717) );
  AOI21XL U7617 ( .A0(n8238), .A1(n3356), .B0(n6351), .Y(n3184) );
  AOI2BB2XL U7618 ( .B0(n6350), .B1(n8224), .A0N(n8224), .A1N(image_data[376]), 
        .Y(n6351) );
  AOI211XL U7619 ( .A0(n3455), .A1(n8114), .B0(n3439), .C0(n6347), .Y(n6350)
         );
  OAI22XL U7620 ( .A0(n3419), .A1(n8381), .B0(n3390), .B1(n6672), .Y(n6347) );
  AOI211XL U7621 ( .A0(n3351), .A1(n8227), .B0(n7175), .C0(n7174), .Y(n3185)
         );
  AOI2BB2XL U7622 ( .B0(n3366), .B1(n8224), .A0N(n8224), .A1N(image_data[377]), 
        .Y(n7174) );
  AOI22XL U7623 ( .A0(n3455), .A1(n7298), .B0(n8238), .B1(n3420), .Y(n7173) );
  AOI211XL U7624 ( .A0(n7795), .A1(n8227), .B0(n7853), .C0(n7852), .Y(n3186)
         );
  AOI2BB2XL U7625 ( .B0(n3348), .B1(n8224), .A0N(n8224), .A1N(image_data[378]), 
        .Y(n7852) );
  AOI22XL U7626 ( .A0(n7923), .A1(n3455), .B0(n8238), .B1(n6880), .Y(n7851) );
  AOI211XL U7627 ( .A0(n3387), .A1(n8227), .B0(n8226), .C0(n8225), .Y(n3187)
         );
  AOI2BB2XL U7628 ( .B0(n3347), .B1(n8224), .A0N(n8224), .A1N(image_data[379]), 
        .Y(n8225) );
  AOI22XL U7629 ( .A0(n3389), .A1(n3455), .B0(n8238), .B1(n6291), .Y(n8223) );
  AOI211XL U7630 ( .A0(n8503), .A1(n8227), .B0(n7413), .C0(n7412), .Y(n3188)
         );
  AOI2BB2XL U7631 ( .B0(n6855), .B1(n8224), .A0N(n8224), .A1N(image_data[380]), 
        .Y(n7412) );
  AOI22XL U7632 ( .A0(n3371), .A1(n3455), .B0(n8238), .B1(n7326), .Y(n7411) );
  AOI211XL U7633 ( .A0(n3361), .A1(n8227), .B0(n7166), .C0(n7165), .Y(n3189)
         );
  AOI2BB2XL U7634 ( .B0(n8496), .B1(n8224), .A0N(n8224), .A1N(image_data[381]), 
        .Y(n7165) );
  AOI22XL U7635 ( .A0(n3357), .A1(n3455), .B0(n8238), .B1(n7078), .Y(n7164) );
  AOI211XL U7636 ( .A0(n3352), .A1(n8227), .B0(n7667), .C0(n7666), .Y(n3190)
         );
  AOI2BB2XL U7637 ( .B0(n3345), .B1(n8224), .A0N(n8224), .A1N(image_data[382]), 
        .Y(n7666) );
  AOI22XL U7638 ( .A0(n3455), .A1(n3353), .B0(n8238), .B1(n3350), .Y(n7665) );
  AOI211XL U7639 ( .A0(n3362), .A1(n8227), .B0(n6676), .C0(n6675), .Y(n3191)
         );
  AOI2BB2XL U7640 ( .B0(n6959), .B1(n8224), .A0N(n8224), .A1N(image_data[383]), 
        .Y(n6675) );
  AOI22XL U7641 ( .A0(n3354), .A1(n3455), .B0(n8238), .B1(n6651), .Y(n6674) );
  AOI21XL U7642 ( .A0(n3373), .A1(n8243), .B0(n6155), .Y(n3192) );
  AOI22XL U7643 ( .A0(n8114), .A1(n8238), .B0(n8378), .B1(n3360), .Y(n6152) );
  AOI211XL U7644 ( .A0(n3351), .A1(n8243), .B0(n7172), .C0(n7171), .Y(n3193)
         );
  AOI2BB2XL U7645 ( .B0(n3366), .B1(n8240), .A0N(n8240), .A1N(image_data[385]), 
        .Y(n7171) );
  AOI22XL U7646 ( .A0(n8238), .A1(n7298), .B0(n8215), .B1(n6332), .Y(n7170) );
  AOI211XL U7647 ( .A0(n7795), .A1(n8243), .B0(n7844), .C0(n7843), .Y(n3194)
         );
  AOI2BB2XL U7648 ( .B0(n3348), .B1(n8240), .A0N(n8240), .A1N(image_data[386]), 
        .Y(n7843) );
  AOI22XL U7649 ( .A0(n7923), .A1(n8238), .B0(n8215), .B1(n6880), .Y(n7842) );
  AOI211XL U7650 ( .A0(n3387), .A1(n8243), .B0(n8242), .C0(n8241), .Y(n3195)
         );
  AOI2BB2XL U7651 ( .B0(n3347), .B1(n8240), .A0N(n8240), .A1N(image_data[387]), 
        .Y(n8241) );
  AOI22XL U7652 ( .A0(n3389), .A1(n8238), .B0(n8378), .B1(n3349), .Y(n8239) );
  AOI21XL U7653 ( .A0(n8503), .A1(n8243), .B0(n6309), .Y(n3196) );
  AOI2BB2XL U7654 ( .B0(n6308), .B1(n8240), .A0N(n8240), .A1N(image_data[388]), 
        .Y(n6309) );
  AOI211XL U7655 ( .A0(n8238), .A1(n3371), .B0(n3418), .C0(n6307), .Y(n6308)
         );
  OAI22XL U7656 ( .A0(n3370), .A1(n8076), .B0(n8055), .B1(n8310), .Y(n6307) );
  AOI211XL U7657 ( .A0(n3361), .A1(n8243), .B0(n7160), .C0(n7159), .Y(n3197)
         );
  AOI2BB2XL U7658 ( .B0(n7303), .B1(n8240), .A0N(n8240), .A1N(image_data[389]), 
        .Y(n7159) );
  AOI22XL U7659 ( .A0(n8378), .A1(n6979), .B0(n8215), .B1(n7078), .Y(n7158) );
  AOI211XL U7660 ( .A0(n3352), .A1(n8243), .B0(n7673), .C0(n7672), .Y(n3198)
         );
  AOI2BB2XL U7661 ( .B0(n3345), .B1(n8240), .A0N(n8240), .A1N(image_data[390]), 
        .Y(n7672) );
  AOI22XL U7662 ( .A0(n8238), .A1(n3353), .B0(n8215), .B1(n3350), .Y(n7671) );
  AOI211XL U7663 ( .A0(n3362), .A1(n8243), .B0(n6664), .C0(n6663), .Y(n3199)
         );
  AOI2BB2XL U7664 ( .B0(n6959), .B1(n8240), .A0N(n8240), .A1N(image_data[391]), 
        .Y(n6663) );
  AOI22XL U7665 ( .A0(n3354), .A1(n8238), .B0(n8215), .B1(n6651), .Y(n6662) );
  AOI211XL U7666 ( .A0(n3373), .A1(n8221), .B0(n7383), .C0(n7382), .Y(n3200)
         );
  AOI2BB2XL U7667 ( .B0(n3344), .B1(n8218), .A0N(n8218), .A1N(image_data[392]), 
        .Y(n7382) );
  AOI22XL U7668 ( .A0(n8114), .A1(n8215), .B0(n8343), .B1(n3360), .Y(n7381) );
  AOI211XL U7669 ( .A0(n3351), .A1(n8221), .B0(n7163), .C0(n7162), .Y(n3201)
         );
  AOI2BB2XL U7670 ( .B0(n3366), .B1(n8218), .A0N(n8218), .A1N(image_data[393]), 
        .Y(n7162) );
  AOI22XL U7671 ( .A0(n8215), .A1(n7298), .B0(n8214), .B1(n6943), .Y(n7161) );
  AOI211XL U7672 ( .A0(n7795), .A1(n8221), .B0(n7832), .C0(n7831), .Y(n3202)
         );
  AOI2BB2XL U7673 ( .B0(n3348), .B1(n8218), .A0N(n8218), .A1N(image_data[394]), 
        .Y(n7831) );
  AOI22XL U7674 ( .A0(n7923), .A1(n8215), .B0(n8214), .B1(n6880), .Y(n7830) );
  AOI211XL U7675 ( .A0(n3387), .A1(n8221), .B0(n8220), .C0(n8219), .Y(n3203)
         );
  AOI2BB2XL U7676 ( .B0(n3347), .B1(n8218), .A0N(n8218), .A1N(image_data[395]), 
        .Y(n8219) );
  AOI22XL U7677 ( .A0(n3389), .A1(n8215), .B0(n8214), .B1(n6291), .Y(n8216) );
  AOI211XL U7678 ( .A0(n8503), .A1(n8221), .B0(n7386), .C0(n7385), .Y(n3204)
         );
  AOI2BB2XL U7679 ( .B0(n6855), .B1(n8218), .A0N(n8218), .A1N(image_data[396]), 
        .Y(n7385) );
  AOI22XL U7680 ( .A0(n3371), .A1(n8215), .B0(n8214), .B1(n7326), .Y(n7384) );
  AOI211XL U7681 ( .A0(n3361), .A1(n8221), .B0(n7127), .C0(n7126), .Y(n3205)
         );
  AOI2BB2XL U7682 ( .B0(n7303), .B1(n8218), .A0N(n8218), .A1N(image_data[397]), 
        .Y(n7126) );
  AOI22XL U7683 ( .A0(n3357), .A1(n8215), .B0(n8214), .B1(n7078), .Y(n7125) );
  AOI211XL U7684 ( .A0(n3352), .A1(n8221), .B0(n7652), .C0(n7651), .Y(n3206)
         );
  AOI2BB2XL U7685 ( .B0(n3345), .B1(n8218), .A0N(n8218), .A1N(image_data[398]), 
        .Y(n7651) );
  AOI22XL U7686 ( .A0(n8343), .A1(n7581), .B0(n8214), .B1(n3350), .Y(n7650) );
  AOI211XL U7687 ( .A0(n3362), .A1(n8221), .B0(n6654), .C0(n6653), .Y(n3207)
         );
  AOI2BB2XL U7688 ( .B0(n6959), .B1(n8218), .A0N(n8218), .A1N(image_data[399]), 
        .Y(n6653) );
  AOI22XL U7689 ( .A0(n8214), .A1(n6651), .B0(n8343), .B1(n3368), .Y(n6652) );
  AOI211XL U7690 ( .A0(n3373), .A1(n8233), .B0(n7389), .C0(n7388), .Y(n3208)
         );
  AOI2BB2XL U7691 ( .B0(n3344), .B1(n8230), .A0N(n8230), .A1N(image_data[400]), 
        .Y(n7388) );
  AOI22XL U7692 ( .A0(n8214), .A1(n8114), .B0(n8228), .B1(n3356), .Y(n7387) );
  AOI211XL U7693 ( .A0(n3351), .A1(n8233), .B0(n7178), .C0(n7177), .Y(n3209)
         );
  AOI2BB2XL U7694 ( .B0(n3366), .B1(n8230), .A0N(n8230), .A1N(image_data[401]), 
        .Y(n7177) );
  AOI22XL U7695 ( .A0(n8214), .A1(n7298), .B0(n8228), .B1(n3420), .Y(n7176) );
  AOI211XL U7696 ( .A0(n7795), .A1(n8233), .B0(n7847), .C0(n7846), .Y(n3210)
         );
  AOI2BB2XL U7697 ( .B0(n3348), .B1(n8230), .A0N(n8230), .A1N(image_data[402]), 
        .Y(n7846) );
  AOI22XL U7698 ( .A0(n7923), .A1(n8214), .B0(n8228), .B1(n7902), .Y(n7845) );
  AOI211XL U7699 ( .A0(n3387), .A1(n8233), .B0(n8232), .C0(n8231), .Y(n3211)
         );
  AOI2BB2XL U7700 ( .B0(n3347), .B1(n8230), .A0N(n8230), .A1N(image_data[403]), 
        .Y(n8231) );
  AOI22XL U7701 ( .A0(n8228), .A1(n6291), .B0(n8342), .B1(n3349), .Y(n8229) );
  AOI211XL U7702 ( .A0(n8503), .A1(n8233), .B0(n7416), .C0(n7415), .Y(n3212)
         );
  AOI2BB2XL U7703 ( .B0(n6855), .B1(n8230), .A0N(n8230), .A1N(image_data[404]), 
        .Y(n7415) );
  AOI22XL U7704 ( .A0(n3371), .A1(n8214), .B0(n8342), .B1(n3388), .Y(n7414) );
  AOI211XL U7705 ( .A0(n3361), .A1(n8233), .B0(n7154), .C0(n7153), .Y(n3213)
         );
  AOI2BB2XL U7706 ( .B0(n7303), .B1(n8230), .A0N(n8230), .A1N(image_data[405]), 
        .Y(n7153) );
  AOI22XL U7707 ( .A0(n7938), .A1(n8214), .B0(n8342), .B1(n6979), .Y(n7152) );
  AOI211XL U7708 ( .A0(n3352), .A1(n8233), .B0(n7676), .C0(n7675), .Y(n3214)
         );
  AOI2BB2XL U7709 ( .B0(n3345), .B1(n8230), .A0N(n8230), .A1N(image_data[406]), 
        .Y(n7675) );
  AOI22XL U7710 ( .A0(n8214), .A1(n3353), .B0(n8228), .B1(n3350), .Y(n7674) );
  AOI211XL U7711 ( .A0(n3362), .A1(n8233), .B0(n6661), .C0(n6660), .Y(n3215)
         );
  AOI2BB2XL U7712 ( .B0(n6959), .B1(n8230), .A0N(n8230), .A1N(image_data[407]), 
        .Y(n6660) );
  AOI22XL U7713 ( .A0(n3354), .A1(n8214), .B0(n8228), .B1(n6651), .Y(n6659) );
  AOI211XL U7714 ( .A0(n3373), .A1(n7352), .B0(n7347), .C0(n7346), .Y(n3216)
         );
  AOI2BB2XL U7715 ( .B0(n3344), .B1(n7349), .A0N(n7349), .A1N(image_data[408]), 
        .Y(n7346) );
  AOI22XL U7716 ( .A0(n8228), .A1(n8114), .B0(n3452), .B1(n3356), .Y(n7345) );
  AOI21XL U7717 ( .A0(n3452), .A1(n6332), .B0(n6335), .Y(n3217) );
  AOI2BB2XL U7718 ( .B0(n6334), .B1(n7349), .A0N(n7349), .A1N(image_data[409]), 
        .Y(n6335) );
  AOI211XL U7719 ( .A0(n8228), .A1(n7298), .B0(n3437), .C0(n6333), .Y(n6334)
         );
  OAI22XL U7720 ( .A0(n3359), .A1(n8329), .B0(n7980), .B1(n6369), .Y(n6333) );
  AOI21XL U7721 ( .A0(n7795), .A1(n7352), .B0(n6286), .Y(n3218) );
  AOI22XL U7722 ( .A0(n7923), .A1(n8228), .B0(n3452), .B1(n7902), .Y(n6283) );
  AOI21XL U7723 ( .A0(n8295), .A1(n3349), .B0(n6372), .Y(n3219) );
  AOI2BB2XL U7724 ( .B0(n6371), .B1(n7349), .A0N(n7349), .A1N(image_data[411]), 
        .Y(n6372) );
  AOI211XL U7725 ( .A0(n8228), .A1(n3389), .B0(n6403), .C0(n6370), .Y(n6371)
         );
  OAI22XL U7726 ( .A0(n8447), .A1(n7864), .B0(n8372), .B1(n6369), .Y(n6370) );
  AOI211XL U7727 ( .A0(n8503), .A1(n7352), .B0(n7351), .C0(n7350), .Y(n3220)
         );
  AOI2BB2XL U7728 ( .B0(n6855), .B1(n7349), .A0N(n7349), .A1N(image_data[412]), 
        .Y(n7350) );
  AOI22XL U7729 ( .A0(n3371), .A1(n8228), .B0(n3452), .B1(n7326), .Y(n7348) );
  AOI211XL U7730 ( .A0(n3361), .A1(n7352), .B0(n7087), .C0(n7086), .Y(n3221)
         );
  AOI2BB2XL U7731 ( .B0(n8496), .B1(n7349), .A0N(n7349), .A1N(image_data[413]), 
        .Y(n7086) );
  AOI22XL U7732 ( .A0(n3357), .A1(n8228), .B0(n8295), .B1(n7261), .Y(n7085) );
  AOI21XL U7733 ( .A0(n3452), .A1(n3350), .B0(n6361), .Y(n3222) );
  AOI2BB2XL U7734 ( .B0(n6360), .B1(n7349), .A0N(n7349), .A1N(image_data[414]), 
        .Y(n6361) );
  AOI211XL U7735 ( .A0(n8295), .A1(n7581), .B0(n3440), .C0(n6359), .Y(n6360)
         );
  OAI22XL U7736 ( .A0(n8509), .A1(n6369), .B0(n3392), .B1(n8159), .Y(n6359) );
  AOI211XL U7737 ( .A0(n3362), .A1(n7352), .B0(n6607), .C0(n6606), .Y(n3223)
         );
  AOI2BB2XL U7738 ( .B0(n6959), .B1(n7349), .A0N(n7349), .A1N(image_data[415]), 
        .Y(n6606) );
  AOI22XL U7739 ( .A0(n3354), .A1(n8228), .B0(n3452), .B1(n6651), .Y(n6605) );
  AOI2BB2XL U7740 ( .B0(n3344), .B1(n8283), .A0N(n8283), .A1N(image_data[416]), 
        .Y(n7456) );
  AOI22XL U7741 ( .A0(n3452), .A1(n8114), .B0(n8492), .B1(n3356), .Y(n7454) );
  AOI211XL U7742 ( .A0(n3351), .A1(n8286), .B0(n7194), .C0(n7193), .Y(n3225)
         );
  AOI2BB2XL U7743 ( .B0(n3366), .B1(n8283), .A0N(n8283), .A1N(image_data[417]), 
        .Y(n7193) );
  AOI22XL U7744 ( .A0(n8294), .A1(n3375), .B0(n8492), .B1(n6332), .Y(n7192) );
  AOI211XL U7745 ( .A0(n7795), .A1(n8286), .B0(n7866), .C0(n7865), .Y(n3226)
         );
  AOI2BB2XL U7746 ( .B0(n3348), .B1(n8283), .A0N(n8283), .A1N(image_data[418]), 
        .Y(n7865) );
  AOI22XL U7747 ( .A0(n8492), .A1(n6880), .B0(n8294), .B1(n3395), .Y(n7863) );
  AOI211XL U7748 ( .A0(n8340), .A1(n8286), .B0(n8285), .C0(n8284), .Y(n3227)
         );
  AOI2BB2XL U7749 ( .B0(n3347), .B1(n8283), .A0N(n8283), .A1N(image_data[419]), 
        .Y(n8284) );
  AOI22XL U7750 ( .A0(n3389), .A1(n3452), .B0(n8294), .B1(n3349), .Y(n8281) );
  AOI2BB2XL U7751 ( .B0(n6855), .B1(n8283), .A0N(n8283), .A1N(image_data[420]), 
        .Y(n7442) );
  AOI22XL U7752 ( .A0(n3371), .A1(n3452), .B0(n8492), .B1(n7326), .Y(n7441) );
  AOI211XL U7753 ( .A0(n3361), .A1(n8286), .B0(n7209), .C0(n7208), .Y(n3229)
         );
  AOI2BB2XL U7754 ( .B0(n8496), .B1(n8283), .A0N(n8283), .A1N(image_data[421]), 
        .Y(n7208) );
  AOI22XL U7755 ( .A0(n3357), .A1(n3452), .B0(n8294), .B1(n7261), .Y(n7207) );
  AOI211XL U7756 ( .A0(n3352), .A1(n8286), .B0(n7693), .C0(n7692), .Y(n3230)
         );
  AOI2BB2XL U7757 ( .B0(n3345), .B1(n8283), .A0N(n8283), .A1N(image_data[422]), 
        .Y(n7692) );
  AOI22XL U7758 ( .A0(n3452), .A1(n3353), .B0(n8294), .B1(n7690), .Y(n7691) );
  AOI211XL U7759 ( .A0(n3362), .A1(n8286), .B0(n6703), .C0(n6702), .Y(n3231)
         );
  AOI2BB2XL U7760 ( .B0(n6959), .B1(n8283), .A0N(n8283), .A1N(image_data[423]), 
        .Y(n6702) );
  AOI22XL U7761 ( .A0(n6973), .A1(n3452), .B0(n8492), .B1(n6651), .Y(n6700) );
  AOI211XL U7762 ( .A0(n3373), .A1(n8128), .B0(n7319), .C0(n7318), .Y(n3232)
         );
  AOI2BB2XL U7763 ( .B0(n3344), .B1(n8498), .A0N(n8498), .A1N(image_data[424]), 
        .Y(n7318) );
  AOI22XL U7764 ( .A0(n8492), .A1(n8114), .B0(n8490), .B1(n3356), .Y(n7316) );
  AOI21XL U7765 ( .A0(n7298), .A1(n8492), .B0(n6331), .Y(n3233) );
  AOI2BB2XL U7766 ( .B0(n6330), .B1(n8498), .A0N(n8498), .A1N(image_data[425]), 
        .Y(n6331) );
  AOI211XL U7767 ( .A0(n3351), .A1(n8493), .B0(n3437), .C0(n6329), .Y(n6330)
         );
  OAI22XL U7768 ( .A0(n3421), .A1(n8125), .B0(n3359), .B1(n7317), .Y(n6329) );
  AOI21XL U7769 ( .A0(n3358), .A1(n8492), .B0(n6380), .Y(n3234) );
  AOI2BB2XL U7770 ( .B0(n6379), .B1(n8498), .A0N(n8498), .A1N(image_data[426]), 
        .Y(n6380) );
  AOI211XL U7771 ( .A0(n8493), .A1(n7795), .B0(n6827), .C0(n6378), .Y(n6379)
         );
  OAI22XL U7772 ( .A0(n3372), .A1(n7317), .B0(n7895), .B1(n8125), .Y(n6378) );
  AOI211XL U7773 ( .A0(n3387), .A1(n8128), .B0(n8127), .C0(n8126), .Y(n3235)
         );
  AOI2BB2XL U7774 ( .B0(n3347), .B1(n8498), .A0N(n8498), .A1N(image_data[427]), 
        .Y(n8126) );
  AOI22XL U7775 ( .A0(n3451), .A1(n3349), .B0(n3389), .B1(n8492), .Y(n8124) );
  AOI211XL U7776 ( .A0(n8503), .A1(n8128), .B0(n7315), .C0(n7314), .Y(n3236)
         );
  AOI2BB2XL U7777 ( .B0(n6855), .B1(n8498), .A0N(n8498), .A1N(image_data[428]), 
        .Y(n7314) );
  AOI22XL U7778 ( .A0(n3451), .A1(n3388), .B0(n8490), .B1(n7487), .Y(n7313) );
  NAND4XL U7779 ( .A(n8496), .B(n8495), .C(n8494), .D(n8498), .Y(n8497) );
  AOI22XL U7780 ( .A0(n3361), .A1(n8493), .B0(n3357), .B1(n8492), .Y(n8494) );
  AOI22XL U7781 ( .A0(n3451), .A1(n6979), .B0(n8490), .B1(n7078), .Y(n8495) );
  AOI211XL U7782 ( .A0(n3352), .A1(n8128), .B0(n7625), .C0(n7624), .Y(n3238)
         );
  AOI2BB2XL U7783 ( .B0(n3345), .B1(n8498), .A0N(n8498), .A1N(image_data[430]), 
        .Y(n7624) );
  AOI22XL U7784 ( .A0(n3451), .A1(n7581), .B0(n8490), .B1(n3350), .Y(n7623) );
  AOI211XL U7785 ( .A0(n6963), .A1(image_data[431]), .B0(n6962), .C0(n6961), 
        .Y(n3239) );
  OAI22XL U7786 ( .A0(n3394), .A1(n7317), .B0(n7578), .B1(n7312), .Y(n6961) );
  AOI21XL U7787 ( .A0(n6959), .A1(n6960), .B0(n6963), .Y(n6962) );
  AOI22XL U7788 ( .A0(n3354), .A1(n8492), .B0(n8490), .B1(n6651), .Y(n6960) );
  AOI2BB2XL U7789 ( .B0(n3344), .B1(n8336), .A0N(n8336), .A1N(image_data[432]), 
        .Y(n7511) );
  AOI22XL U7790 ( .A0(n8490), .A1(n8114), .B0(n7513), .B1(n3356), .Y(n7510) );
  AOI211XL U7791 ( .A0(n3351), .A1(n8339), .B0(n6942), .C0(n6941), .Y(n3241)
         );
  AOI2BB2XL U7792 ( .B0(n3346), .B1(n8336), .A0N(n8336), .A1N(image_data[433]), 
        .Y(n6941) );
  AOI22XL U7793 ( .A0(n8490), .A1(n7298), .B0(n7513), .B1(n6332), .Y(n6940) );
  AOI211XL U7794 ( .A0(n7795), .A1(n8339), .B0(n7897), .C0(n7896), .Y(n3242)
         );
  AOI2BB2XL U7795 ( .B0(n3348), .B1(n8336), .A0N(n8336), .A1N(image_data[434]), 
        .Y(n7896) );
  AOI22XL U7796 ( .A0(n8334), .A1(n7761), .B0(n3358), .B1(n8490), .Y(n7894) );
  AOI211XL U7797 ( .A0(n8340), .A1(n8339), .B0(n8338), .C0(n8337), .Y(n3243)
         );
  AOI2BB2XL U7798 ( .B0(n3347), .B1(n8336), .A0N(n8336), .A1N(image_data[435]), 
        .Y(n8337) );
  AOI22XL U7799 ( .A0(n8334), .A1(n3349), .B0(n3389), .B1(n8490), .Y(n8335) );
  AOI2BB2XL U7800 ( .B0(n6855), .B1(n8336), .A0N(n8336), .A1N(image_data[436]), 
        .Y(n7515) );
  AOI22XL U7801 ( .A0(n8334), .A1(n3388), .B0(n7513), .B1(n7326), .Y(n7514) );
  AOI211XL U7802 ( .A0(n3361), .A1(n8339), .B0(n6851), .C0(n6850), .Y(n3245)
         );
  AOI2BB2XL U7803 ( .B0(n8496), .B1(n8336), .A0N(n8336), .A1N(image_data[437]), 
        .Y(n6850) );
  AOI22XL U7804 ( .A0(n7938), .A1(n8490), .B0(n7513), .B1(n7078), .Y(n6849) );
  AOI211XL U7805 ( .A0(n3352), .A1(n8339), .B0(n7722), .C0(n7721), .Y(n3246)
         );
  AOI2BB2XL U7806 ( .B0(n3345), .B1(n8336), .A0N(n8336), .A1N(image_data[438]), 
        .Y(n7721) );
  AOI22XL U7807 ( .A0(n8334), .A1(n7581), .B0(n3353), .B1(n8490), .Y(n7720) );
  AOI211XL U7808 ( .A0(n3362), .A1(n8339), .B0(n6746), .C0(n6745), .Y(n3247)
         );
  AOI2BB2XL U7809 ( .B0(n6586), .B1(n8336), .A0N(n8336), .A1N(image_data[439]), 
        .Y(n6745) );
  AOI22XL U7810 ( .A0(n6973), .A1(n8490), .B0(n8334), .B1(n3368), .Y(n6743) );
  AOI211XL U7811 ( .A0(n3373), .A1(n8384), .B0(n7493), .C0(n7492), .Y(n3248)
         );
  AOI2BB2XL U7812 ( .B0(n3344), .B1(n7874), .A0N(n7874), .A1N(image_data[440]), 
        .Y(n7492) );
  AOI22XL U7813 ( .A0(n8377), .A1(n3360), .B0(n8378), .B1(n3356), .Y(n7491) );
  AOI211XL U7814 ( .A0(n3351), .A1(n8384), .B0(n6927), .C0(n6926), .Y(n3249)
         );
  AOI2BB2XL U7815 ( .B0(n3346), .B1(n7874), .A0N(n7874), .A1N(image_data[441]), 
        .Y(n6926) );
  AOI22XL U7816 ( .A0(n8377), .A1(n3375), .B0(n8378), .B1(n6332), .Y(n6925) );
  AOI211XL U7817 ( .A0(n7795), .A1(n8384), .B0(n7876), .C0(n7875), .Y(n3250)
         );
  AOI2BB2XL U7818 ( .B0(n3348), .B1(n7874), .A0N(n7874), .A1N(image_data[442]), 
        .Y(n7875) );
  AOI22XL U7819 ( .A0(n8378), .A1(n6880), .B0(n8377), .B1(n3395), .Y(n7873) );
  AOI211XL U7820 ( .A0(n8384), .A1(n3369), .B0(n8383), .C0(n8382), .Y(n3251)
         );
  OAI2BB2XL U7821 ( .B0(n6407), .B1(n8381), .A0N(n8380), .A1N(image_data[443]), 
        .Y(n8382) );
  AOI21XL U7822 ( .A0(n3347), .A1(n8379), .B0(n8380), .Y(n8383) );
  AOI22XL U7823 ( .A0(n8378), .A1(n6291), .B0(n8377), .B1(n8376), .Y(n8379) );
  AOI211XL U7824 ( .A0(n8503), .A1(n8384), .B0(n7490), .C0(n7489), .Y(n3252)
         );
  AOI2BB2XL U7825 ( .B0(n6855), .B1(n7874), .A0N(n7874), .A1N(image_data[444]), 
        .Y(n7489) );
  AOI22XL U7826 ( .A0(n8377), .A1(n3388), .B0(n8378), .B1(n7487), .Y(n7488) );
  AOI211XL U7827 ( .A0(n3361), .A1(n8384), .B0(n7245), .C0(n7244), .Y(n3253)
         );
  AOI2BB2XL U7828 ( .B0(n7303), .B1(n7874), .A0N(n7874), .A1N(image_data[445]), 
        .Y(n7244) );
  AOI22XL U7829 ( .A0(n8377), .A1(n6979), .B0(n8378), .B1(n7078), .Y(n7243) );
  AOI211XL U7830 ( .A0(n3352), .A1(n8384), .B0(n7707), .C0(n7706), .Y(n3254)
         );
  AOI2BB2XL U7831 ( .B0(n3345), .B1(n7874), .A0N(n7874), .A1N(image_data[446]), 
        .Y(n7706) );
  AOI22XL U7832 ( .A0(n8377), .A1(n7581), .B0(n8378), .B1(n3350), .Y(n7705) );
  AOI211XL U7833 ( .A0(n3362), .A1(n8384), .B0(n6908), .C0(n6907), .Y(n3255)
         );
  AOI2BB2XL U7834 ( .B0(n6959), .B1(n7874), .A0N(n7874), .A1N(image_data[447]), 
        .Y(n6907) );
  AOI22XL U7835 ( .A0(n8378), .A1(n6651), .B0(n8377), .B1(n3368), .Y(n6906) );
  OAI22XL U7836 ( .A0(n3419), .A1(n8323), .B0(n8111), .B1(n8076), .Y(n8077) );
  AOI22XL U7837 ( .A0(n3373), .A1(n8074), .B0(n8343), .B1(n3356), .Y(n8075) );
  AOI211XL U7838 ( .A0(n3351), .A1(n3436), .B0(n6930), .C0(n6929), .Y(n3257)
         );
  AOI2BB2XL U7839 ( .B0(n3346), .B1(n8324), .A0N(n8324), .A1N(image_data[449]), 
        .Y(n6929) );
  AOI22XL U7840 ( .A0(n8378), .A1(n7298), .B0(n8343), .B1(n6943), .Y(n6928) );
  AOI211XL U7841 ( .A0(n7795), .A1(n3436), .B0(n7886), .C0(n7885), .Y(n3258)
         );
  AOI2BB2XL U7842 ( .B0(n3348), .B1(n8324), .A0N(n8324), .A1N(image_data[450]), 
        .Y(n7885) );
  AOI22XL U7843 ( .A0(n7923), .A1(n8378), .B0(n8343), .B1(n6880), .Y(n7884) );
  AOI211XL U7844 ( .A0(n3387), .A1(n3436), .B0(n8326), .C0(n8325), .Y(n3259)
         );
  AOI2BB2XL U7845 ( .B0(n3347), .B1(n8324), .A0N(n8324), .A1N(image_data[451]), 
        .Y(n8325) );
  AOI22XL U7846 ( .A0(n3389), .A1(n8378), .B0(n8343), .B1(n8341), .Y(n8322) );
  AOI21XL U7847 ( .A0(n8503), .A1(n3436), .B0(n6135), .Y(n3260) );
  AOI22XL U7848 ( .A0(n8438), .A1(n3388), .B0(n3371), .B1(n8378), .Y(n6133) );
  AOI211XL U7849 ( .A0(n3436), .A1(n3361), .B0(n7933), .C0(n7932), .Y(n3261)
         );
  OAI2BB2XL U7850 ( .B0(n3391), .B1(n8076), .A0N(n8079), .A1N(image_data[453]), 
        .Y(n7932) );
  AOI22XL U7851 ( .A0(n8438), .A1(n6979), .B0(n8343), .B1(n7930), .Y(n7931) );
  AOI211XL U7852 ( .A0(n3352), .A1(n3436), .B0(n7713), .C0(n7712), .Y(n3262)
         );
  AOI2BB2XL U7853 ( .B0(n3345), .B1(n8324), .A0N(n8324), .A1N(image_data[454]), 
        .Y(n7712) );
  AOI22XL U7854 ( .A0(n8438), .A1(n7581), .B0(n3353), .B1(n8378), .Y(n7711) );
  AOI211XL U7855 ( .A0(n3362), .A1(n3436), .B0(n6911), .C0(n6910), .Y(n3263)
         );
  AOI2BB2XL U7856 ( .B0(n6959), .B1(n8324), .A0N(n8324), .A1N(image_data[455]), 
        .Y(n6910) );
  AOI22XL U7857 ( .A0(n6973), .A1(n8378), .B0(n8343), .B1(n6651), .Y(n6909) );
  AOI2BB2XL U7858 ( .B0(n3344), .B1(n8345), .A0N(n8345), .A1N(image_data[456]), 
        .Y(n7519) );
  AOI22XL U7859 ( .A0(n8343), .A1(n8114), .B0(n8342), .B1(n7517), .Y(n7518) );
  AOI211XL U7860 ( .A0(n3351), .A1(n8348), .B0(n6946), .C0(n6945), .Y(n3265)
         );
  AOI2BB2XL U7861 ( .B0(n3346), .B1(n8345), .A0N(n8345), .A1N(image_data[457]), 
        .Y(n6945) );
  AOI22XL U7862 ( .A0(n8343), .A1(n7298), .B0(n8342), .B1(n6943), .Y(n6944) );
  AOI211XL U7863 ( .A0(n7795), .A1(n8348), .B0(n7905), .C0(n7904), .Y(n3266)
         );
  AOI2BB2XL U7864 ( .B0(n3348), .B1(n8345), .A0N(n8345), .A1N(image_data[458]), 
        .Y(n7904) );
  AOI22XL U7865 ( .A0(n3358), .A1(n8343), .B0(n8342), .B1(n7902), .Y(n7903) );
  AOI211XL U7866 ( .A0(n3387), .A1(n8348), .B0(n8347), .C0(n8346), .Y(n3267)
         );
  AOI2BB2XL U7867 ( .B0(n3347), .B1(n8345), .A0N(n8345), .A1N(image_data[459]), 
        .Y(n8346) );
  AOI22XL U7868 ( .A0(n3389), .A1(n8343), .B0(n8342), .B1(n8341), .Y(n8344) );
  AOI211XL U7869 ( .A0(n8503), .A1(n8348), .B0(n6877), .C0(n6876), .Y(n3268)
         );
  AOI2BB2XL U7870 ( .B0(n6855), .B1(n8345), .A0N(n8345), .A1N(image_data[460]), 
        .Y(n6876) );
  AOI22XL U7871 ( .A0(n3371), .A1(n8343), .B0(n8342), .B1(n7487), .Y(n6874) );
  AOI211XL U7872 ( .A0(n3361), .A1(n8348), .B0(n7264), .C0(n7263), .Y(n3269)
         );
  AOI2BB2XL U7873 ( .B0(n8496), .B1(n8345), .A0N(n8345), .A1N(image_data[461]), 
        .Y(n7263) );
  AOI22XL U7874 ( .A0(n3357), .A1(n8343), .B0(n8182), .B1(n7261), .Y(n7262) );
  AOI2BB2XL U7875 ( .B0(n3345), .B1(n8345), .A0N(n8345), .A1N(image_data[462]), 
        .Y(n7725) );
  AOI22XL U7876 ( .A0(n8343), .A1(n3353), .B0(n8342), .B1(n7723), .Y(n7724) );
  AOI211XL U7877 ( .A0(n3362), .A1(n8348), .B0(n6917), .C0(n6916), .Y(n3271)
         );
  AOI2BB2XL U7878 ( .B0(n6959), .B1(n8345), .A0N(n8345), .A1N(image_data[463]), 
        .Y(n6916) );
  AOI22XL U7879 ( .A0(n3354), .A1(n8343), .B0(n8342), .B1(n6651), .Y(n6915) );
  AOI2BB2XL U7880 ( .B0(n3367), .B1(n8330), .A0N(n8330), .A1N(image_data[464]), 
        .Y(n6814) );
  AOI22XL U7881 ( .A0(n8114), .A1(n8342), .B0(n8513), .B1(n3360), .Y(n6813) );
  AOI2BB2XL U7882 ( .B0(n3346), .B1(n8330), .A0N(n8330), .A1N(image_data[465]), 
        .Y(n6932) );
  AOI22XL U7883 ( .A0(n7298), .A1(n8342), .B0(n8513), .B1(n3375), .Y(n6931) );
  AOI22XL U7884 ( .A0(n3358), .A1(n8342), .B0(n8295), .B1(n7902), .Y(n5600) );
  AOI2BB2XL U7885 ( .B0(n3347), .B1(n8330), .A0N(n8330), .A1N(image_data[467]), 
        .Y(n8331) );
  AOI22XL U7886 ( .A0(n3389), .A1(n8342), .B0(n8513), .B1(n8376), .Y(n8328) );
  AOI2BB2XL U7887 ( .B0(n6855), .B1(n8330), .A0N(n8330), .A1N(image_data[468]), 
        .Y(n6865) );
  AOI22XL U7888 ( .A0(n3371), .A1(n8342), .B0(n8513), .B1(n3388), .Y(n6864) );
  AOI221XL U7889 ( .A0(image_data[469]), .A1(n7311), .B0(n7310), .B1(n8330), 
        .C0(n7309), .Y(n3277) );
  AOI22XL U7890 ( .A0(n8513), .A1(n6979), .B0(n8295), .B1(n7930), .Y(n7308) );
  NOR2XL U7891 ( .A(n3396), .B(n8329), .Y(n6887) );
  AOI32XL U7892 ( .A0(n3365), .A1(n8330), .A2(n6885), .B0(n7311), .B1(n8553), 
        .Y(n6886) );
  AOI22XL U7893 ( .A0(n8342), .A1(n6951), .B0(n8513), .B1(n7690), .Y(n6885) );
  AOI2BB2XL U7894 ( .B0(n6959), .B1(n8330), .A0N(n8330), .A1N(image_data[471]), 
        .Y(n6913) );
  AOI22XL U7895 ( .A0(n3354), .A1(n8342), .B0(n8513), .B1(n3368), .Y(n6912) );
  AOI211XL U7896 ( .A0(n3373), .A1(n8300), .B0(n6818), .C0(n6817), .Y(n3280)
         );
  AOI2BB2XL U7897 ( .B0(n3367), .B1(n8297), .A0N(n8297), .A1N(image_data[472]), 
        .Y(n6817) );
  AOI22XL U7898 ( .A0(n8295), .A1(n8114), .B0(n8294), .B1(n7517), .Y(n6816) );
  AOI211XL U7899 ( .A0(n3351), .A1(n8300), .B0(n6939), .C0(n6938), .Y(n3281)
         );
  AOI2BB2XL U7900 ( .B0(n3346), .B1(n8297), .A0N(n8297), .A1N(image_data[473]), 
        .Y(n6938) );
  AOI22XL U7901 ( .A0(n8295), .A1(n7298), .B0(n8294), .B1(n6943), .Y(n6937) );
  AOI211XL U7902 ( .A0(n7795), .A1(n8300), .B0(n6835), .C0(n6834), .Y(n3282)
         );
  AOI2BB2XL U7903 ( .B0(n3348), .B1(n8297), .A0N(n8297), .A1N(image_data[474]), 
        .Y(n6834) );
  AOI22XL U7904 ( .A0(n3358), .A1(n8295), .B0(n8294), .B1(n7902), .Y(n6833) );
  AOI211XL U7905 ( .A0(n3369), .A1(n8300), .B0(n8299), .C0(n8298), .Y(n3283)
         );
  AOI2BB2XL U7906 ( .B0(n3347), .B1(n8297), .A0N(n8297), .A1N(image_data[475]), 
        .Y(n8298) );
  AOI22XL U7907 ( .A0(n8423), .A1(n8295), .B0(n8294), .B1(n8341), .Y(n8296) );
  AOI211XL U7908 ( .A0(n8503), .A1(n8300), .B0(n6869), .C0(n6868), .Y(n3284)
         );
  AOI2BB2XL U7909 ( .B0(n6855), .B1(n8297), .A0N(n8297), .A1N(image_data[476]), 
        .Y(n6868) );
  AOI22XL U7910 ( .A0(n7377), .A1(n8295), .B0(n8294), .B1(n7487), .Y(n6867) );
  AOI211XL U7911 ( .A0(n3361), .A1(n8300), .B0(n6848), .C0(n6847), .Y(n3285)
         );
  AOI2BB2XL U7912 ( .B0(n8496), .B1(n8297), .A0N(n8297), .A1N(image_data[477]), 
        .Y(n6847) );
  AOI22XL U7913 ( .A0(n3357), .A1(n8295), .B0(n8294), .B1(n7930), .Y(n6846) );
  AOI211XL U7914 ( .A0(n3352), .A1(n8300), .B0(n6808), .C0(n6807), .Y(n3286)
         );
  AOI2BB2XL U7915 ( .B0(n3365), .B1(n8297), .A0N(n8297), .A1N(image_data[478]), 
        .Y(n6807) );
  AOI22XL U7916 ( .A0(n8295), .A1(n3353), .B0(n8294), .B1(n7723), .Y(n6805) );
  AOI211XL U7917 ( .A0(n3362), .A1(n8300), .B0(n6901), .C0(n6900), .Y(n3287)
         );
  AOI2BB2XL U7918 ( .B0(n6959), .B1(n8297), .A0N(n8297), .A1N(image_data[479]), 
        .Y(n6900) );
  AOI22XL U7919 ( .A0(n6973), .A1(n8295), .B0(n8294), .B1(n6651), .Y(n6899) );
  AOI211XL U7920 ( .A0(n3373), .A1(n8253), .B0(n6812), .C0(n6811), .Y(n3288)
         );
  AOI2BB2XL U7921 ( .B0(n3367), .B1(n8250), .A0N(n8250), .A1N(image_data[480]), 
        .Y(n6811) );
  AOI22XL U7922 ( .A0(n3451), .A1(n3356), .B0(n8114), .B1(n8294), .Y(n6809) );
  AOI211XL U7923 ( .A0(n3351), .A1(n8253), .B0(n6921), .C0(n6920), .Y(n3289)
         );
  AOI2BB2XL U7924 ( .B0(n3346), .B1(n8250), .A0N(n8250), .A1N(image_data[481]), 
        .Y(n6920) );
  AOI22XL U7925 ( .A0(n3451), .A1(n6332), .B0(n7298), .B1(n8294), .Y(n6918) );
  AOI211XL U7926 ( .A0(n7795), .A1(n8253), .B0(n7850), .C0(n7849), .Y(n3290)
         );
  AOI2BB2XL U7927 ( .B0(n3348), .B1(n8250), .A0N(n8250), .A1N(image_data[482]), 
        .Y(n7849) );
  AOI22XL U7928 ( .A0(n3451), .A1(n6880), .B0(n3358), .B1(n8294), .Y(n7848) );
  AOI211XL U7929 ( .A0(n8340), .A1(n8253), .B0(n8252), .C0(n8251), .Y(n3291)
         );
  AOI2BB2XL U7930 ( .B0(n3347), .B1(n8250), .A0N(n8250), .A1N(image_data[483]), 
        .Y(n8251) );
  AOI22XL U7931 ( .A0(n3451), .A1(n6291), .B0(n8423), .B1(n8294), .Y(n8249) );
  AOI211XL U7932 ( .A0(n8503), .A1(n8253), .B0(n6860), .C0(n6859), .Y(n3292)
         );
  AOI2BB2XL U7933 ( .B0(n6855), .B1(n8250), .A0N(n8250), .A1N(image_data[484]), 
        .Y(n6859) );
  AOI22XL U7934 ( .A0(n3451), .A1(n7326), .B0(n3371), .B1(n8294), .Y(n6858) );
  AOI211XL U7935 ( .A0(n3361), .A1(n8253), .B0(n6839), .C0(n6838), .Y(n3293)
         );
  AOI2BB2XL U7936 ( .B0(n7303), .B1(n8250), .A0N(n8250), .A1N(image_data[485]), 
        .Y(n6838) );
  AOI22XL U7937 ( .A0(n3451), .A1(n7078), .B0(n3357), .B1(n8294), .Y(n6836) );
  AOI211XL U7938 ( .A0(n3352), .A1(n8253), .B0(n6799), .C0(n6798), .Y(n3294)
         );
  AOI2BB2XL U7939 ( .B0(n3365), .B1(n8250), .A0N(n8250), .A1N(image_data[486]), 
        .Y(n6798) );
  AOI22XL U7940 ( .A0(n3451), .A1(n3350), .B0(n6951), .B1(n8294), .Y(n6796) );
  AOI211XL U7941 ( .A0(n3362), .A1(n8253), .B0(n6895), .C0(n6894), .Y(n3295)
         );
  AOI2BB2XL U7942 ( .B0(n6959), .B1(n8250), .A0N(n8250), .A1N(image_data[487]), 
        .Y(n6894) );
  AOI22XL U7943 ( .A0(n6973), .A1(n8294), .B0(n3451), .B1(n7035), .Y(n6892) );
  AOI211XL U7944 ( .A0(n3425), .A1(image_data[488]), .B0(n8072), .C0(n8071), 
        .Y(n3296) );
  OAI22XL U7945 ( .A0(n3385), .A1(n8070), .B0(n8069), .B1(n3390), .Y(n8071) );
  AOI21XL U7946 ( .A0(n3367), .A1(n8068), .B0(n3425), .Y(n8072) );
  AOI22XL U7947 ( .A0(n3376), .A1(n3360), .B0(n3451), .B1(n8114), .Y(n8068) );
  AOI211XL U7948 ( .A0(n3425), .A1(image_data[489]), .B0(n7982), .C0(n7981), 
        .Y(n3297) );
  OAI22XL U7949 ( .A0(n3421), .A1(n8070), .B0(n8069), .B1(n7980), .Y(n7981) );
  AOI21XL U7950 ( .A0(n3366), .A1(n7979), .B0(n3425), .Y(n7982) );
  AOI22XL U7951 ( .A0(n3376), .A1(n3375), .B0(n3451), .B1(n7298), .Y(n7979) );
  AOI211XL U7952 ( .A0(n6891), .A1(n7795), .B0(n6832), .C0(n6831), .Y(n3298)
         );
  AOI2BB2XL U7953 ( .B0(n3348), .B1(n6957), .A0N(n6957), .A1N(image_data[490]), 
        .Y(n6831) );
  AOI22XL U7954 ( .A0(n3376), .A1(n7761), .B0(n3451), .B1(n3358), .Y(n6830) );
  AOI211XL U7955 ( .A0(n6891), .A1(n3369), .B0(n6405), .C0(n6404), .Y(n3299)
         );
  AOI2BB2XL U7956 ( .B0(n3347), .B1(n6957), .A0N(n6957), .A1N(image_data[491]), 
        .Y(n6404) );
  AOI22XL U7957 ( .A0(n3376), .A1(n3349), .B0(n3451), .B1(n8423), .Y(n6402) );
  AOI211XL U7958 ( .A0(n6891), .A1(n8503), .B0(n6863), .C0(n6862), .Y(n3300)
         );
  AOI2BB2XL U7959 ( .B0(n6855), .B1(n6957), .A0N(n6957), .A1N(image_data[492]), 
        .Y(n6862) );
  AOI22XL U7960 ( .A0(n3376), .A1(n3388), .B0(n3451), .B1(n3371), .Y(n6861) );
  AOI211XL U7961 ( .A0(n6891), .A1(n3361), .B0(n6845), .C0(n6844), .Y(n3301)
         );
  AOI2BB2XL U7962 ( .B0(n8496), .B1(n6957), .A0N(n6957), .A1N(image_data[493]), 
        .Y(n6844) );
  AOI22XL U7963 ( .A0(n3376), .A1(n6979), .B0(n3451), .B1(n3357), .Y(n6843) );
  AOI221XL U7964 ( .A0(image_data[494]), .A1(n3425), .B0(n6958), .B1(n6957), 
        .C0(n6956), .Y(n3302) );
  AOI22XL U7965 ( .A0(n3376), .A1(n7581), .B0(n3451), .B1(n3353), .Y(n6955) );
  AOI211XL U7966 ( .A0(n3362), .A1(n6891), .B0(n6890), .C0(n6889), .Y(n3303)
         );
  AOI2BB2XL U7967 ( .B0(n6959), .B1(n6957), .A0N(n6957), .A1N(image_data[495]), 
        .Y(n6889) );
  AOI22XL U7968 ( .A0(n3376), .A1(n3368), .B0(n3354), .B1(n3451), .Y(n6888) );
  AOI211XL U7969 ( .A0(n3373), .A1(n8248), .B0(n7422), .C0(n7421), .Y(n3304)
         );
  AOI2BB2XL U7970 ( .B0(n3344), .B1(n8245), .A0N(n8245), .A1N(image_data[496]), 
        .Y(n7421) );
  AOI22XL U7971 ( .A0(n8334), .A1(n8114), .B0(n8377), .B1(n3356), .Y(n7420) );
  AOI211XL U7972 ( .A0(n3351), .A1(n8248), .B0(n6924), .C0(n6923), .Y(n3305)
         );
  AOI2BB2XL U7973 ( .B0(n3346), .B1(n8245), .A0N(n8245), .A1N(image_data[497]), 
        .Y(n6923) );
  AOI22XL U7974 ( .A0(n8334), .A1(n7298), .B0(n8377), .B1(n6332), .Y(n6922) );
  AOI211XL U7975 ( .A0(n7795), .A1(n8248), .B0(n6829), .C0(n6828), .Y(n3306)
         );
  AOI2BB2XL U7976 ( .B0(n3348), .B1(n8245), .A0N(n8245), .A1N(image_data[498]), 
        .Y(n6828) );
  AOI22XL U7977 ( .A0(n8334), .A1(n3358), .B0(n8377), .B1(n6880), .Y(n6826) );
  AOI211XL U7978 ( .A0(n8340), .A1(n8248), .B0(n8247), .C0(n8246), .Y(n3307)
         );
  AOI2BB2XL U7979 ( .B0(n3347), .B1(n8245), .A0N(n8245), .A1N(image_data[499]), 
        .Y(n8246) );
  AOI22XL U7980 ( .A0(n8334), .A1(n3389), .B0(n8377), .B1(n8341), .Y(n8244) );
  AOI211XL U7981 ( .A0(n8503), .A1(n8248), .B0(n6857), .C0(n6856), .Y(n3308)
         );
  AOI2BB2XL U7982 ( .B0(n6855), .B1(n8245), .A0N(n8245), .A1N(image_data[500]), 
        .Y(n6856) );
  AOI22XL U7983 ( .A0(n8334), .A1(n3371), .B0(n8377), .B1(n7326), .Y(n6853) );
  AOI211XL U7984 ( .A0(n3361), .A1(n8248), .B0(n6842), .C0(n6841), .Y(n3309)
         );
  AOI2BB2XL U7985 ( .B0(n8496), .B1(n8245), .A0N(n8245), .A1N(image_data[501]), 
        .Y(n6841) );
  AOI22XL U7986 ( .A0(n8334), .A1(n3357), .B0(n8377), .B1(n7078), .Y(n6840) );
  AOI211XL U7987 ( .A0(n3352), .A1(n8248), .B0(n7670), .C0(n7669), .Y(n3310)
         );
  AOI2BB2XL U7988 ( .B0(n3345), .B1(n8245), .A0N(n8245), .A1N(image_data[502]), 
        .Y(n7669) );
  AOI22XL U7989 ( .A0(n8334), .A1(n3353), .B0(n8377), .B1(n3350), .Y(n7668) );
  AOI211XL U7990 ( .A0(n3362), .A1(n8248), .B0(n6898), .C0(n6897), .Y(n3311)
         );
  AOI2BB2XL U7991 ( .B0(n6959), .B1(n8245), .A0N(n8245), .A1N(image_data[503]), 
        .Y(n6897) );
  AOI22XL U7992 ( .A0(n6973), .A1(n8334), .B0(n8377), .B1(n7035), .Y(n6896) );
  AOI211XL U7993 ( .A0(n3355), .A1(n8444), .B0(n8120), .C0(n8119), .Y(n3312)
         );
  AOI2BB2XL U7994 ( .B0(n3367), .B1(n8441), .A0N(n8441), .A1N(image_data[504]), 
        .Y(n8119) );
  AOI22XL U7995 ( .A0(n8114), .A1(n8377), .B0(n8437), .B1(n3360), .Y(n8118) );
  AOI211XL U7996 ( .A0(n3351), .A1(n8444), .B0(n8012), .C0(n8011), .Y(n3313)
         );
  AOI2BB2XL U7997 ( .B0(n3346), .B1(n8441), .A0N(n8441), .A1N(image_data[505]), 
        .Y(n8011) );
  AOI22XL U7998 ( .A0(n7298), .A1(n8377), .B0(n8437), .B1(n3375), .Y(n8010) );
  AOI211XL U7999 ( .A0(n7795), .A1(n8444), .B0(n7788), .C0(n7787), .Y(n3314)
         );
  AOI2BB2XL U8000 ( .B0(n3348), .B1(n8441), .A0N(n8441), .A1N(image_data[506]), 
        .Y(n7787) );
  AOI22XL U8001 ( .A0(n3358), .A1(n8377), .B0(n8437), .B1(n3395), .Y(n7786) );
  AOI211XL U8002 ( .A0(n3369), .A1(n8444), .B0(n8443), .C0(n8442), .Y(n3315)
         );
  AOI2BB2XL U8003 ( .B0(n3347), .B1(n8441), .A0N(n8441), .A1N(image_data[507]), 
        .Y(n8442) );
  AOI22XL U8004 ( .A0(n8438), .A1(n6291), .B0(n8437), .B1(n3349), .Y(n8439) );
  AOI211XL U8005 ( .A0(n8503), .A1(n8444), .B0(n8067), .C0(n8066), .Y(n3316)
         );
  AOI2BB2XL U8006 ( .B0(n6855), .B1(n8441), .A0N(n8441), .A1N(image_data[508]), 
        .Y(n8066) );
  AOI22XL U8007 ( .A0(n8438), .A1(n7326), .B0(n3371), .B1(n8377), .Y(n8065) );
  AOI211XL U8008 ( .A0(n3361), .A1(n8444), .B0(n7968), .C0(n7967), .Y(n3317)
         );
  AOI2BB2XL U8009 ( .B0(n8496), .B1(n8441), .A0N(n8441), .A1N(image_data[509]), 
        .Y(n7967) );
  AOI22XL U8010 ( .A0(n8438), .A1(n7078), .B0(n8437), .B1(n6979), .Y(n7966) );
  AOI211XL U8011 ( .A0(n3352), .A1(n8444), .B0(n7618), .C0(n7617), .Y(n3318)
         );
  AOI2BB2XL U8012 ( .B0(n3365), .B1(n8441), .A0N(n8441), .A1N(image_data[510]), 
        .Y(n7617) );
  AOI22XL U8013 ( .A0(n8377), .A1(n3353), .B0(n8437), .B1(n7581), .Y(n7616) );
  AOI211XL U8014 ( .A0(n3362), .A1(n8444), .B0(n7048), .C0(n7047), .Y(n3319)
         );
  AOI2BB2XL U8015 ( .B0(n6959), .B1(n8441), .A0N(n8441), .A1N(image_data[511]), 
        .Y(n7047) );
  AOI22XL U8016 ( .A0(n3354), .A1(n8377), .B0(n8437), .B1(n3368), .Y(n7045) );
  AOI211XL U8017 ( .A0(op4[4]), .A1(n6321), .B0(n6385), .C0(n6320), .Y(n3325)
         );
  AOI211XL U8018 ( .A0(n6319), .A1(n6318), .B0(op4[4]), .C0(n6317), .Y(n6320)
         );
  AOI22XL U8019 ( .A0(cmd_valid), .A1(cmd[0]), .B0(cmd_reg[0]), .B1(n6388), 
        .Y(n3334) );
  AOI22XL U8020 ( .A0(cmd_valid), .A1(cmd[1]), .B0(cmd_reg[1]), .B1(n6388), 
        .Y(n3335) );
  AOI22XL U8021 ( .A0(cmd_valid), .A1(cmd[2]), .B0(cmd_reg[2]), .B1(n6388), 
        .Y(n3336) );
  AOI22XL U8022 ( .A0(cmd_valid), .A1(cmd[3]), .B0(cmd_reg[3]), .B1(n6388), 
        .Y(n3337) );
  NAND2X2 U8023 ( .A(n6825), .B(n6646), .Y(n3405) );
  OR3XL U8024 ( .A(n6721), .B(n8302), .C(n6723), .Y(n3406) );
  OR3XL U8025 ( .A(n8452), .B(n7023), .C(n7021), .Y(n3407) );
  OR3XL U8026 ( .A(n3384), .B(n6770), .C(n7014), .Y(n3408) );
  OR3XL U8027 ( .A(n8315), .B(n6643), .C(n6640), .Y(n3409) );
  NOR4X2 U8028 ( .A(n4584), .B(n4583), .C(n4582), .D(n4581), .Y(n4585) );
  NOR4X2 U8029 ( .A(n5312), .B(n5311), .C(n5310), .D(n5309), .Y(n5313) );
  NOR4X2 U8030 ( .A(n5354), .B(n5353), .C(n5352), .D(n5351), .Y(n5355) );
  NOR4X2 U8031 ( .A(n5396), .B(n5395), .C(n5394), .D(n5393), .Y(n5397) );
  NOR4X2 U8032 ( .A(n5438), .B(n5437), .C(n5436), .D(n5435), .Y(n5439) );
  NOR4X2 U8033 ( .A(n5480), .B(n5479), .C(n5478), .D(n5477), .Y(n5481) );
  NOR4X2 U8034 ( .A(n5522), .B(n5521), .C(n5520), .D(n5519), .Y(n5523) );
  NOR4X2 U8035 ( .A(n5596), .B(n5595), .C(n5594), .D(n5593), .Y(n5597) );
  NOR4X2 U8036 ( .A(n4564), .B(n4563), .C(n4562), .D(n4561), .Y(n4586) );
  NOR4X2 U8037 ( .A(n5292), .B(n5291), .C(n5290), .D(n5289), .Y(n5314) );
  NOR4X2 U8038 ( .A(n5334), .B(n5333), .C(n5332), .D(n5331), .Y(n5356) );
  NOR4X2 U8039 ( .A(n5376), .B(n5375), .C(n5374), .D(n5373), .Y(n5398) );
  NOR4X2 U8040 ( .A(n5418), .B(n5417), .C(n5416), .D(n5415), .Y(n5440) );
  NOR4X2 U8041 ( .A(n5460), .B(n5459), .C(n5458), .D(n5457), .Y(n5482) );
  NOR4X2 U8042 ( .A(n5502), .B(n5501), .C(n5500), .D(n5499), .Y(n5524) );
  NOR4X2 U8043 ( .A(n5544), .B(n5543), .C(n5542), .D(n5541), .Y(n5598) );
  NOR2X4 U8044 ( .A(n8521), .B(n8489), .Y(IRAM_A[5]) );
  NOR2X4 U8045 ( .A(n8520), .B(n8489), .Y(IRAM_A[1]) );
  AOI22X2 U8046 ( .A0(n4871), .A1(n6421), .B0(n8459), .B1(n6420), .Y(n7068) );
  NAND2X1 U8047 ( .A(n8467), .B(n6639), .Y(n8202) );
  INVXL U8048 ( .A(n7058), .Y(n3411) );
  INVX1 U8049 ( .A(N2772), .Y(n5115) );
  INVX1 U8050 ( .A(n8500), .Y(n3413) );
  AOI21XL U8051 ( .A0(n6760), .A1(n7031), .B0(n6159), .Y(n6163) );
  AOI21XL U8052 ( .A0(n6688), .A1(n6760), .B0(n6687), .Y(n6691) );
  INVXL U8053 ( .A(n8375), .Y(n3414) );
  INVX1 U8054 ( .A(n3414), .Y(n3415) );
  AOI21XL U8055 ( .A0(n7032), .A1(n6871), .B0(n5930), .Y(n8375) );
  AOI21XL U8056 ( .A0(n6986), .A1(n6688), .B0(n6666), .Y(n6667) );
  AOI21XL U8057 ( .A0(n6986), .A1(n7031), .B0(n6614), .Y(n6615) );
  AOI21XL U8058 ( .A0(n6904), .A1(n7031), .B0(n6656), .Y(n6657) );
  AOI21XL U8059 ( .A0(n6904), .A1(n6688), .B0(n6150), .Y(n6154) );
  INVXL U8060 ( .A(n8517), .Y(n3416) );
  INVX1 U8061 ( .A(n3416), .Y(n3417) );
  OAI21XL U8062 ( .A0(n5799), .A1(n6583), .B0(n5798), .Y(n6854) );
  NAND2X1 U8063 ( .A(op4[3]), .B(n6984), .Y(n6710) );
  INVXL U8064 ( .A(n8014), .Y(n3420) );
  CLKINVX3 U8065 ( .A(n3420), .Y(n3421) );
  INVXL U8066 ( .A(n6968), .Y(n3422) );
  INVX1 U8067 ( .A(n3422), .Y(n3423) );
  AOI21XL U8068 ( .A0(n6994), .A1(n6779), .B0(n6390), .Y(n6968) );
  INVXL U8069 ( .A(n8073), .Y(n3424) );
  INVX1 U8070 ( .A(n3424), .Y(n3425) );
  AOI21XL U8071 ( .A0(n6872), .A1(n6779), .B0(n6399), .Y(n8073) );
  AOI21XL U8072 ( .A0(n8496), .A1(n7931), .B0(n8079), .Y(n7933) );
  AOI21XL U8073 ( .A0(n3367), .A1(n8075), .B0(n8079), .Y(n8078) );
  OAI221XL U8074 ( .A0(n8079), .A1(n6134), .B0(n8324), .B1(n8557), .C0(n6133), 
        .Y(n6135) );
  NAND2X4 U8075 ( .A(n4535), .B(n8527), .Y(n4549) );
  CLKINVX3 U8076 ( .A(n3404), .Y(n3430) );
  NOR2X4 U8077 ( .A(n8526), .B(n8489), .Y(IRAM_A[0]) );
  NOR2X2 U8078 ( .A(n3438), .B(n6902), .Y(n6742) );
  INVX4 U8079 ( .A(reset), .Y(n8578) );
  INVX4 U8080 ( .A(reset), .Y(n8577) );
  INVX4 U8081 ( .A(reset), .Y(n8576) );
  INVX4 U8082 ( .A(reset), .Y(n8583) );
  INVX4 U8083 ( .A(reset), .Y(n8579) );
  INVX4 U8084 ( .A(reset), .Y(n8595) );
  NOR2X2 U8085 ( .A(n8524), .B(n7033), .Y(n5929) );
  NOR2X2 U8086 ( .A(n8524), .B(n6902), .Y(n6825) );
  NAND2X2 U8087 ( .A(op4[4]), .B(op4[5]), .Y(n6902) );
  CLKINVX3 U8088 ( .A(n3401), .Y(n3432) );
  INVXL U8089 ( .A(n8272), .Y(n3433) );
  INVXL U8090 ( .A(n8327), .Y(n3435) );
  OAI21XL U8091 ( .A0(n5697), .A1(n6583), .B0(n5696), .Y(n6919) );
  NOR2X2 U8092 ( .A(n6287), .B(n7039), .Y(n6872) );
  NOR2X2 U8093 ( .A(n6673), .B(n6672), .Y(n8227) );
  NOR2X2 U8094 ( .A(n6678), .B(n6677), .Y(n8258) );
  AOI21XL U8095 ( .A0(n6994), .A1(n6688), .B0(n6343), .Y(n6678) );
  NOR2X2 U8096 ( .A(n6683), .B(n6682), .Y(n8265) );
  NAND2X2 U8097 ( .A(n8480), .B(n8527), .Y(n6275) );
  OAI221XL U8098 ( .A0(in_valid), .A1(IRAM_D[4]), .B0(n8523), .B1(IROM_Q[4]), 
        .C0(n8480), .Y(n5798) );
  OAI221XL U8099 ( .A0(in_valid), .A1(IRAM_D[5]), .B0(n8523), .B1(IROM_Q[5]), 
        .C0(n8480), .Y(n6019) );
  OAI221XL U8100 ( .A0(in_valid), .A1(IRAM_D[6]), .B0(n8523), .B1(IROM_Q[6]), 
        .C0(n8480), .Y(n5901) );
  NOR2X4 U8101 ( .A(cs[0]), .B(cs[1]), .Y(n8480) );
  NAND2X4 U8102 ( .A(op2[0]), .B(op2[1]), .Y(n4588) );
  OAI21XL U8103 ( .A0(n6122), .A1(n6583), .B0(n6121), .Y(n6810) );
  OAI21XL U8104 ( .A0(n5902), .A1(n6583), .B0(n5901), .Y(n6797) );
  NAND2X4 U8105 ( .A(n6820), .B(n6992), .Y(n8419) );
  CLKINVX2 U8106 ( .A(n8483), .Y(n6992) );
  NOR2X4 U8107 ( .A(n5013), .B(op4[5]), .Y(n6820) );
  CLKINVX3 U8108 ( .A(n3403), .Y(n3443) );
  CLKINVX3 U8109 ( .A(n3403), .Y(n3444) );
  CLKINVX3 U8110 ( .A(n3402), .Y(n3445) );
  CLKINVX3 U8111 ( .A(n3402), .Y(n3446) );
  BUFX1 U8112 ( .A(n6750), .Y(n3449) );
  NAND2X2 U8113 ( .A(n6647), .B(n3449), .Y(n6650) );
  NAND2X2 U8114 ( .A(n6820), .B(n3449), .Y(n8370) );
  NAND2X2 U8115 ( .A(n6646), .B(n5929), .Y(n8101) );
  NOR2X4 U8116 ( .A(n5002), .B(op2[2]), .Y(n8467) );
  NAND2X2 U8117 ( .A(n6136), .B(op4[5]), .Y(n6728) );
  NAND2X2 U8118 ( .A(n8524), .B(n6721), .Y(n8304) );
  NAND3X2 U8119 ( .A(n8529), .B(n8528), .C(op2[1]), .Y(n7034) );
  INVX4 U8120 ( .A(reset), .Y(n8571) );
  OAI21XL U8121 ( .A0(n6136), .A1(n8525), .B0(n6802), .Y(n5167) );
  NOR2X4 U8122 ( .A(n8524), .B(n6665), .Y(n8141) );
  NAND2X4 U8123 ( .A(n6984), .B(n8524), .Y(n6766) );
  NOR2X4 U8124 ( .A(n8518), .B(op4[5]), .Y(n6984) );
  NAND2X4 U8125 ( .A(n6820), .B(n6699), .Y(n8446) );
  NOR2X4 U8126 ( .A(n8527), .B(n8489), .Y(IRAM_A[4]) );
  NOR2X4 U8127 ( .A(n8522), .B(n8489), .Y(IRAM_A[3]) );
  NAND2X4 U8128 ( .A(cs[0]), .B(cs[1]), .Y(n8489) );
  AOI21X1 U8129 ( .A0(n6904), .A1(n7040), .B0(n6903), .Y(n8380) );
  INVX12 U8130 ( .A(n3374), .Y(n7298) );
  INVXL U8131 ( .A(n7029), .Y(n3453) );
  NOR2X2 U8132 ( .A(n5928), .B(n6583), .Y(n7938) );
  CLKINVX3 U8133 ( .A(n7377), .Y(n8035) );
  NOR2X1 U8134 ( .A(n3482), .B(n3476), .Y(n4713) );
  NAND2X2 U8135 ( .A(n6030), .B(n6646), .Y(n8267) );
  NOR2X2 U8136 ( .A(n7564), .B(n7560), .Y(n8429) );
  AOI21XL U8137 ( .A0(n6879), .A1(n8333), .B0(n5602), .Y(n3274) );
  NOR2X2 U8138 ( .A(n7003), .B(n7002), .Y(n7769) );
  NOR2X2 U8139 ( .A(n3417), .B(n8508), .Y(n8416) );
  AOI21XL U8140 ( .A0(n7032), .A1(n7031), .B0(n7030), .Y(n8517) );
  AOI221X4 U8141 ( .A0(n6415), .A1(n5705), .B0(n6416), .B1(n5704), .C0(n6027), 
        .Y(n8503) );
  NAND2X2 U8142 ( .A(n6384), .B(n6304), .Y(n6416) );
  CLKINVX2 U8143 ( .A(n8079), .Y(n8324) );
  INVXL U8144 ( .A(n8018), .Y(n3454) );
  AOI21XL U8145 ( .A0(n6855), .A1(n8027), .B0(n3454), .Y(n8030) );
  AOI21XL U8146 ( .A0(n3365), .A1(n7583), .B0(n3454), .Y(n7585) );
  AOI21XL U8147 ( .A0(n7096), .A1(n6871), .B0(n6366), .Y(n8028) );
  NAND2X4 U8148 ( .A(n8526), .B(n8520), .Y(n3461) );
  NAND2X2 U8149 ( .A(n8526), .B(n8520), .Y(n4536) );
  NAND2X4 U8150 ( .A(n3449), .B(n6142), .Y(n8351) );
  CLKINVX2 U8151 ( .A(n3415), .Y(n8096) );
  AOI21XL U8152 ( .A0(n8021), .A1(n8165), .B0(n3363), .Y(n6993) );
  NAND2X2 U8153 ( .A(n6151), .B(n6647), .Y(n8165) );
  NAND2X1 U8154 ( .A(op4[3]), .B(n6620), .Y(n8184) );
  INVX1 U8155 ( .A(n4868), .Y(n3465) );
  NOR2X2 U8156 ( .A(n6777), .B(n6728), .Y(n7826) );
  NAND3X4 U8157 ( .A(n8530), .B(op2[0]), .C(op2[2]), .Y(n6777) );
  AOI22X4 U8158 ( .A0(IROM_A[5]), .A1(n5482), .B0(n5481), .B1(n8521), .Y(
        IRAM_D[4]) );
  CLKINVX2 U8159 ( .A(n7973), .Y(n7980) );
  OAI21XL U8160 ( .A0(n5094), .A1(n5093), .B0(n5092), .Y(n5095) );
  AOI21XL U8161 ( .A0(n5142), .A1(n4991), .B0(n5140), .Y(n4994) );
  AOI21XL U8162 ( .A0(n6634), .A1(n6631), .B0(n3363), .Y(n6632) );
  AOI21XL U8163 ( .A0(n6650), .A1(n6658), .B0(n3363), .Y(n6648) );
  AOI21XL U8164 ( .A0(n6992), .A1(n6984), .B0(n8273), .Y(n6987) );
  AOI21XL U8165 ( .A0(n5910), .A1(n7864), .B0(n3363), .Y(n5909) );
  AOI21XL U8166 ( .A0(n7008), .A1(n6872), .B0(n6793), .Y(n6794) );
  AOI21XL U8167 ( .A0(n7096), .A1(n7095), .B0(n7094), .Y(n7575) );
  AOI21XL U8168 ( .A0(n8503), .A1(n8397), .B0(n5805), .Y(n2932) );
  AOI21XL U8169 ( .A0(n3369), .A1(n7922), .B0(n6295), .Y(n2987) );
  NOR2X1 U8170 ( .A(op2[1]), .B(op2[0]), .Y(n5809) );
  CLKINVX3 U8171 ( .A(n5809), .Y(n5002) );
  NOR2X2 U8172 ( .A(n6401), .B(op4[4]), .Y(n6136) );
  NAND2X2 U8173 ( .A(n8467), .B(n6136), .Y(n5010) );
  NAND2X2 U8174 ( .A(op4[4]), .B(n3470), .Y(n3482) );
  NAND3X2 U8175 ( .A(n6401), .B(n8518), .C(n8528), .Y(n3483) );
  NOR2X1 U8176 ( .A(n5002), .B(n3483), .Y(n4670) );
  NOR2X1 U8177 ( .A(n5002), .B(n3484), .Y(n4768) );
  NAND3X1 U8178 ( .A(op2[2]), .B(n8518), .C(n8524), .Y(n3485) );
  NOR2X1 U8179 ( .A(n5002), .B(n3485), .Y(n3792) );
  NOR2X4 U8180 ( .A(n5002), .B(n3432), .Y(n4702) );
  NAND3X2 U8181 ( .A(op2[2]), .B(n6401), .C(n8518), .Y(n3486) );
  NOR2X2 U8182 ( .A(n5002), .B(n3486), .Y(n3791) );
  NOR2X1 U8183 ( .A(n3481), .B(n3471), .Y(n3797) );
  NOR2X4 U8184 ( .A(n3482), .B(n3471), .Y(n4707) );
  NOR2X2 U8185 ( .A(n3483), .B(n3471), .Y(n4708) );
  NOR2X1 U8186 ( .A(n3485), .B(n3471), .Y(n3799) );
  NOR2X4 U8187 ( .A(n3432), .B(n3471), .Y(n4763) );
  NAND2X2 U8188 ( .A(op2[0]), .B(n8530), .Y(n3476) );
  NOR2X1 U8189 ( .A(n3481), .B(n3476), .Y(n3804) );
  NOR2X2 U8190 ( .A(n3483), .B(n3476), .Y(n4753) );
  NOR2X1 U8191 ( .A(n3485), .B(n3476), .Y(n3805) );
  NOR2X4 U8192 ( .A(n3432), .B(n3476), .Y(n4714) );
  NOR2X2 U8193 ( .A(n3486), .B(n3476), .Y(n4754) );
  NOR2X1 U8194 ( .A(n3481), .B(n4588), .Y(n3810) );
  NOR2X4 U8195 ( .A(n3482), .B(n4588), .Y(n4719) );
  NOR2X2 U8196 ( .A(n3483), .B(n4588), .Y(n4720) );
  NOR2X1 U8197 ( .A(n3485), .B(n4588), .Y(n3811) );
  NOR2X4 U8198 ( .A(n3432), .B(n4588), .Y(n4721) );
  NOR2X2 U8199 ( .A(n3486), .B(n4588), .Y(n4722) );
  NAND2X1 U8200 ( .A(n8467), .B(n6353), .Y(n7041) );
  NOR2X4 U8201 ( .A(n7041), .B(n6401), .Y(n8438) );
  OAI2BB1X4 U8202 ( .A0N(op4[5]), .A1N(n5010), .B0(n8323), .Y(n5165) );
  AOI22X2 U8203 ( .A0(n5165), .A1(n3685), .B0(n3684), .B1(n4777), .Y(N2782) );
  AOI22X2 U8204 ( .A0(n3450), .A1(n3770), .B0(n3769), .B1(n4959), .Y(N2759) );
  AOI22X2 U8205 ( .A0(n5165), .A1(n3863), .B0(n3862), .B1(n4777), .Y(N2784) );
  NAND2X2 U8206 ( .A(n6401), .B(n5009), .Y(n6131) );
  NAND2X1 U8207 ( .A(n6131), .B(n8518), .Y(n3864) );
  AOI2BB2X4 U8208 ( .B0(n8525), .B1(n3864), .A0N(n3864), .A1N(n8525), .Y(n5168) );
  NOR4X2 U8209 ( .A(n4000), .B(n3999), .C(n3998), .D(n3997), .Y(n4022) );
  NOR4X2 U8210 ( .A(n4020), .B(n4019), .C(n4018), .D(n4017), .Y(n4021) );
  AOI22X4 U8211 ( .A0(op4[5]), .A1(n4022), .B0(n4021), .B1(n8525), .Y(N2765)
         );
  AOI22X2 U8212 ( .A0(n5165), .A1(n4149), .B0(n4148), .B1(n4777), .Y(N2783) );
  NOR4X2 U8213 ( .A(n4211), .B(n4210), .C(n4209), .D(n4208), .Y(n4233) );
  NOR4X2 U8214 ( .A(n4231), .B(n4230), .C(n4229), .D(n4228), .Y(n4232) );
  AOI22X4 U8215 ( .A0(n5168), .A1(n4233), .B0(n4232), .B1(n4868), .Y(N2773) );
  NOR4X2 U8216 ( .A(n4253), .B(n4252), .C(n4251), .D(n4250), .Y(n4275) );
  NOR4X2 U8217 ( .A(n4273), .B(n4272), .C(n4271), .D(n4270), .Y(n4274) );
  AOI22X4 U8218 ( .A0(n3465), .A1(n4275), .B0(n4274), .B1(n4868), .Y(N2774) );
  NOR4X2 U8219 ( .A(n4295), .B(n4294), .C(n4293), .D(n4292), .Y(n4317) );
  NOR4X2 U8220 ( .A(n4315), .B(n4314), .C(n4313), .D(n4312), .Y(n4316) );
  AOI22X4 U8221 ( .A0(n5168), .A1(n4317), .B0(n4316), .B1(n4868), .Y(N2775) );
  AOI22X2 U8222 ( .A0(n5168), .A1(n4359), .B0(n4358), .B1(n4868), .Y(N2772) );
  AOI22X2 U8223 ( .A0(n3450), .A1(n4534), .B0(n4533), .B1(n4959), .Y(N2757) );
  NOR2X1 U8224 ( .A(IROM_A[2]), .B(IROM_A[3]), .Y(n4535) );
  NOR2X4 U8225 ( .A(n3461), .B(n4549), .Y(n5546) );
  NOR2X4 U8226 ( .A(n3461), .B(n3430), .Y(n5545) );
  NAND3X4 U8227 ( .A(IROM_A[3]), .B(n8527), .C(n8519), .Y(n4550) );
  NOR2X4 U8228 ( .A(n3461), .B(n4550), .Y(n5548) );
  NAND3X4 U8229 ( .A(IROM_A[4]), .B(IROM_A[3]), .C(n8519), .Y(n4551) );
  NOR2X4 U8230 ( .A(n4536), .B(n4551), .Y(n5547) );
  NAND3X4 U8231 ( .A(IROM_A[2]), .B(n8527), .C(n8522), .Y(n4552) );
  NOR2X4 U8232 ( .A(n3461), .B(n4552), .Y(n5550) );
  NAND3X4 U8233 ( .A(IROM_A[2]), .B(IROM_A[4]), .C(n8522), .Y(n4553) );
  NOR2X4 U8234 ( .A(n4536), .B(n4553), .Y(n5549) );
  NAND3X4 U8235 ( .A(IROM_A[2]), .B(IROM_A[3]), .C(n8527), .Y(n4554) );
  NOR2X4 U8236 ( .A(n3461), .B(n4554), .Y(n5552) );
  NAND3X4 U8237 ( .A(IROM_A[4]), .B(IROM_A[2]), .C(IROM_A[3]), .Y(n4556) );
  NOR2X4 U8238 ( .A(n4536), .B(n4556), .Y(n5551) );
  NOR2X4 U8239 ( .A(n4549), .B(n3444), .Y(n5558) );
  NOR2X4 U8240 ( .A(n3430), .B(n3443), .Y(n5557) );
  NOR2X4 U8241 ( .A(n4550), .B(n3444), .Y(n5560) );
  NOR2X4 U8242 ( .A(n4551), .B(n3443), .Y(n5559) );
  NOR2X4 U8243 ( .A(n4552), .B(n3444), .Y(n5562) );
  NOR2X4 U8244 ( .A(n4553), .B(n3443), .Y(n5561) );
  NOR2X4 U8245 ( .A(n4554), .B(n3444), .Y(n5564) );
  NOR2X4 U8246 ( .A(n4556), .B(n3443), .Y(n5563) );
  NOR2X4 U8247 ( .A(n4549), .B(n3446), .Y(n5570) );
  NOR2X4 U8248 ( .A(n3430), .B(n3445), .Y(n5569) );
  NOR2X4 U8249 ( .A(n4550), .B(n3446), .Y(n5572) );
  NOR2X4 U8250 ( .A(n4551), .B(n3445), .Y(n5571) );
  NOR2X4 U8251 ( .A(n4552), .B(n3446), .Y(n5574) );
  NOR2X4 U8252 ( .A(n4553), .B(n3445), .Y(n5573) );
  NOR2X4 U8253 ( .A(n4554), .B(n3446), .Y(n5576) );
  NOR2X4 U8254 ( .A(n4556), .B(n3445), .Y(n5575) );
  NOR2X4 U8255 ( .A(n4549), .B(n3456), .Y(n5582) );
  NOR2X4 U8256 ( .A(n3430), .B(n3456), .Y(n5581) );
  NOR2X4 U8257 ( .A(n4550), .B(n3456), .Y(n5584) );
  NOR2X4 U8258 ( .A(n4551), .B(n3456), .Y(n5583) );
  NOR2X4 U8259 ( .A(n4552), .B(n3456), .Y(n5586) );
  NOR2X4 U8260 ( .A(n4553), .B(n3456), .Y(n5585) );
  NOR2X4 U8261 ( .A(n4554), .B(n3456), .Y(n5588) );
  NOR2X4 U8262 ( .A(n4556), .B(n3456), .Y(n5587) );
  AOI22X4 U8263 ( .A0(IROM_A[5]), .A1(n4586), .B0(n4585), .B1(n8521), .Y(
        IRAM_D[2]) );
  INVX1 U8264 ( .A(n6303), .Y(n6384) );
  CLKINVX2 U8265 ( .A(n6416), .Y(n6415) );
  NAND2X1 U8266 ( .A(n8532), .B(cmd_reg[3]), .Y(n5268) );
  NOR2X2 U8267 ( .A(n5268), .B(n6416), .Y(n6417) );
  NOR2X1 U8268 ( .A(cs[0]), .B(n8533), .Y(n4590) );
  NOR2X1 U8269 ( .A(n6583), .B(n5268), .Y(n6414) );
  OAI21XL U8270 ( .A0(N2784), .A1(n6417), .B0(n6414), .Y(n4587) );
  AOI21XL U8271 ( .A0(n6415), .A1(n4986), .B0(n4587), .Y(n6879) );
  NOR3X2 U8272 ( .A(IROM_A[5]), .B(n8522), .C(n6275), .Y(n7096) );
  NOR3X2 U8273 ( .A(IROM_A[0]), .B(IROM_A[2]), .C(n8520), .Y(n7031) );
  NOR2X1 U8274 ( .A(n8528), .B(n5809), .Y(n5706) );
  CLKINVX3 U8275 ( .A(n6281), .Y(n7029) );
  INVX1 U8276 ( .A(n6353), .Y(n7033) );
  NOR2X4 U8277 ( .A(n7034), .B(n6766), .Y(n8259) );
  NOR2X4 U8278 ( .A(n7029), .B(n6766), .Y(n8404) );
  AOI31X1 U8279 ( .A0(n4595), .A1(n4590), .A2(n6311), .B0(n6414), .Y(n6337) );
  AOI21X1 U8280 ( .A0(n7096), .A1(n7031), .B0(n4591), .Y(n7564) );
  INVX1 U8281 ( .A(n6414), .Y(n6027) );
  BUFX3 U8282 ( .A(n4593), .Y(n6421) );
  BUFX3 U8283 ( .A(n4594), .Y(n6420) );
  INVX1 U8284 ( .A(n7754), .Y(n7761) );
  AOI22X2 U8285 ( .A0(n5165), .A1(n4680), .B0(n4679), .B1(n4777), .Y(n5698) );
  AOI22X2 U8286 ( .A0(op4[5]), .A1(n4732), .B0(n4731), .B1(n8525), .Y(n8459)
         );
  AOI22X2 U8287 ( .A0(n5165), .A1(n4779), .B0(n4778), .B1(n4777), .Y(n6123) );
  OAI21XL U8288 ( .A0(n4780), .A1(n5150), .B0(n5151), .Y(n4781) );
  OAI21XL U8289 ( .A0(n4782), .A1(n5156), .B0(n5155), .Y(n4783) );
  AOI22X2 U8290 ( .A0(n5168), .A1(n4827), .B0(n4826), .B1(n4868), .Y(n6127) );
  OAI21XL U8291 ( .A0(N2775), .A1(n4979), .B0(n4873), .Y(n4874) );
  OAI21XL U8292 ( .A0(n4875), .A1(n5113), .B0(n5112), .Y(n4876) );
  OAI21XL U8293 ( .A0(N2755), .A1(N2779), .B0(n5118), .Y(n4976) );
  AOI22X1 U8294 ( .A0(n3450), .A1(n4918), .B0(n4917), .B1(n4959), .Y(n6124) );
  AOI22X2 U8295 ( .A0(n3450), .A1(n4961), .B0(n4960), .B1(n4959), .Y(n8458) );
  INVX1 U8296 ( .A(n6124), .Y(n6028) );
  OAI21XL U8297 ( .A0(n4980), .A1(n5127), .B0(n5126), .Y(n4982) );
  OAI21XL U8298 ( .A0(n4983), .A1(n5133), .B0(n5132), .Y(n4996) );
  OAI21XL U8299 ( .A0(n4994), .A1(n5144), .B0(n5143), .Y(n4995) );
  NAND2X2 U8300 ( .A(n5001), .B(n5000), .Y(n6498) );
  OAI21X2 U8301 ( .A0(n8530), .A1(n5004), .B0(n5003), .Y(n5042) );
  NOR2X2 U8302 ( .A(n5706), .B(n8467), .Y(n5174) );
  AOI22X4 U8303 ( .A0(n5005), .A1(n8528), .B0(n5174), .B1(n5004), .Y(n5023) );
  OAI21XL U8304 ( .A0(n6401), .A1(n5009), .B0(n6131), .Y(n5178) );
  OAI221X4 U8305 ( .A0(n5180), .A1(n5008), .B0(n5178), .B1(n5007), .C0(n5006), 
        .Y(n5022) );
  NOR2X2 U8306 ( .A(n5023), .B(n5022), .Y(n5018) );
  OAI21XL U8307 ( .A0(n6151), .A1(n8518), .B0(n5010), .Y(n5181) );
  AOI22X1 U8308 ( .A0(n5012), .A1(n5181), .B0(n5011), .B1(op4[4]), .Y(n5017)
         );
  OAI21XL U8309 ( .A0(n8518), .A1(n8524), .B0(n5013), .Y(n5186) );
  AOI22X1 U8310 ( .A0(n5015), .A1(n5184), .B0(n5014), .B1(n5186), .Y(n5016) );
  NAND2X4 U8311 ( .A(n5017), .B(n5016), .Y(n5024) );
  CLKINVX3 U8312 ( .A(n5024), .Y(n5021) );
  NAND2X4 U8313 ( .A(n5018), .B(n5021), .Y(n5044) );
  NOR2X4 U8314 ( .A(n3462), .B(n5044), .Y(n6444) );
  NAND2X4 U8315 ( .A(n5024), .B(n5018), .Y(n5045) );
  NOR2X4 U8316 ( .A(n3462), .B(n5045), .Y(n6443) );
  NAND3X4 U8317 ( .A(n5022), .B(n5021), .C(n5019), .Y(n5046) );
  NOR2X4 U8318 ( .A(n3462), .B(n5046), .Y(n6446) );
  NAND3X4 U8319 ( .A(n5024), .B(n5022), .C(n5019), .Y(n5047) );
  NOR2X4 U8320 ( .A(n3462), .B(n5047), .Y(n6445) );
  NAND3X4 U8321 ( .A(n5023), .B(n5021), .C(n5020), .Y(n5048) );
  NOR2X4 U8322 ( .A(n3462), .B(n5048), .Y(n6448) );
  NAND3X4 U8323 ( .A(n5023), .B(n5024), .C(n5020), .Y(n5049) );
  NOR2X4 U8324 ( .A(n3462), .B(n5049), .Y(n6447) );
  NAND3X4 U8325 ( .A(n5023), .B(n5022), .C(n5021), .Y(n5050) );
  NOR2X4 U8326 ( .A(n3462), .B(n5050), .Y(n6450) );
  NAND3X4 U8327 ( .A(n5024), .B(n5023), .C(n5022), .Y(n5052) );
  NOR2X4 U8328 ( .A(n3462), .B(n5052), .Y(n6449) );
  NAND2X4 U8329 ( .A(n5042), .B(n5030), .Y(n5031) );
  NOR2X4 U8330 ( .A(n5044), .B(n5031), .Y(n6456) );
  NOR2X4 U8331 ( .A(n5045), .B(n5031), .Y(n6455) );
  NOR2X4 U8332 ( .A(n5046), .B(n5031), .Y(n6458) );
  NOR2X4 U8333 ( .A(n5047), .B(n3447), .Y(n6457) );
  NOR2X4 U8334 ( .A(n5048), .B(n5031), .Y(n6460) );
  NOR2X4 U8335 ( .A(n5049), .B(n3447), .Y(n6459) );
  NOR2X4 U8336 ( .A(n5050), .B(n3447), .Y(n6462) );
  NOR2X4 U8337 ( .A(n5052), .B(n3447), .Y(n6461) );
  NOR2X4 U8338 ( .A(n5044), .B(n3458), .Y(n6468) );
  NOR2X4 U8339 ( .A(n5045), .B(n3458), .Y(n6467) );
  NOR2X4 U8340 ( .A(n5046), .B(n3458), .Y(n6470) );
  NOR2X4 U8341 ( .A(n5047), .B(n3458), .Y(n6469) );
  NOR2X4 U8342 ( .A(n5048), .B(n3458), .Y(n6472) );
  NOR2X4 U8343 ( .A(n5049), .B(n3458), .Y(n6471) );
  NOR2X4 U8344 ( .A(n5050), .B(n3458), .Y(n6474) );
  NOR2X4 U8345 ( .A(n5052), .B(n3458), .Y(n6473) );
  NOR2X4 U8346 ( .A(n5044), .B(n3457), .Y(n6480) );
  NOR2X4 U8347 ( .A(n5045), .B(n3457), .Y(n6479) );
  NOR2X4 U8348 ( .A(n5046), .B(n3457), .Y(n6482) );
  NOR2X4 U8349 ( .A(n5047), .B(n3457), .Y(n6481) );
  NOR2X4 U8350 ( .A(n5048), .B(n3457), .Y(n6484) );
  NOR2X4 U8351 ( .A(n5049), .B(n3457), .Y(n6483) );
  NOR2X4 U8352 ( .A(n5050), .B(n3457), .Y(n6486) );
  NOR2X4 U8353 ( .A(n5052), .B(n3457), .Y(n6485) );
  OAI21XL U8354 ( .A0(n5102), .A1(n5101), .B0(n5100), .Y(n5104) );
  OAI21XL U8355 ( .A0(n5114), .A1(n5113), .B0(n5112), .Y(n5116) );
  OAI21XL U8356 ( .A0(n5128), .A1(n5127), .B0(n5126), .Y(n5130) );
  OAI21XL U8357 ( .A0(n5134), .A1(n5133), .B0(n5132), .Y(n5147) );
  OAI21XL U8358 ( .A0(n5139), .A1(n5138), .B0(n5137), .Y(n5141) );
  OAI21XL U8359 ( .A0(n5145), .A1(n5144), .B0(n5143), .Y(n5146) );
  OAI21XL U8360 ( .A0(n5157), .A1(n5156), .B0(n5155), .Y(n5158) );
  NAND2X2 U8361 ( .A(n5170), .B(n5169), .Y(n6574) );
  OAI21X2 U8362 ( .A0(n8530), .A1(n5173), .B0(n5172), .Y(n5214) );
  AOI22X4 U8363 ( .A0(n5175), .A1(n8528), .B0(n5174), .B1(n5173), .Y(n5195) );
  OAI221X4 U8364 ( .A0(n5180), .A1(n5179), .B0(n5178), .B1(n5177), .C0(n5176), 
        .Y(n5194) );
  NOR2X2 U8365 ( .A(n5195), .B(n5194), .Y(n5190) );
  AOI22X1 U8366 ( .A0(op4[4]), .A1(n5183), .B0(n5182), .B1(n5181), .Y(n5189)
         );
  AOI22X1 U8367 ( .A0(n5187), .A1(n5186), .B0(n5185), .B1(n5184), .Y(n5188) );
  NAND2X4 U8368 ( .A(n5189), .B(n5188), .Y(n5196) );
  CLKINVX3 U8369 ( .A(n5196), .Y(n5193) );
  NAND2X4 U8370 ( .A(n5190), .B(n5193), .Y(n5216) );
  NOR2X4 U8371 ( .A(n3463), .B(n5216), .Y(n6520) );
  NAND2X4 U8372 ( .A(n5196), .B(n5190), .Y(n5217) );
  NOR2X4 U8373 ( .A(n3463), .B(n5217), .Y(n6519) );
  NAND3X4 U8374 ( .A(n5194), .B(n5193), .C(n5191), .Y(n5218) );
  NOR2X4 U8375 ( .A(n3463), .B(n5218), .Y(n6522) );
  NAND3X4 U8376 ( .A(n5196), .B(n5194), .C(n5191), .Y(n5219) );
  NOR2X4 U8377 ( .A(n3463), .B(n5219), .Y(n6521) );
  NAND3X4 U8378 ( .A(n5195), .B(n5193), .C(n5192), .Y(n5220) );
  NOR2X4 U8379 ( .A(n3463), .B(n5220), .Y(n6524) );
  NAND3X4 U8380 ( .A(n5195), .B(n5196), .C(n5192), .Y(n5221) );
  NOR2X4 U8381 ( .A(n3463), .B(n5221), .Y(n6523) );
  NAND3X4 U8382 ( .A(n5195), .B(n5194), .C(n5193), .Y(n5222) );
  NOR2X4 U8383 ( .A(n3463), .B(n5222), .Y(n6526) );
  NAND3X4 U8384 ( .A(n5196), .B(n5195), .C(n5194), .Y(n5224) );
  NOR2X4 U8385 ( .A(n3463), .B(n5224), .Y(n6525) );
  NAND2X4 U8386 ( .A(n5214), .B(n5202), .Y(n5203) );
  NOR2X4 U8387 ( .A(n5216), .B(n5203), .Y(n6532) );
  NOR2X4 U8388 ( .A(n5217), .B(n5203), .Y(n6531) );
  NOR2X4 U8389 ( .A(n5218), .B(n5203), .Y(n6534) );
  NOR2X4 U8390 ( .A(n5219), .B(n3448), .Y(n6533) );
  NOR2X4 U8391 ( .A(n5220), .B(n5203), .Y(n6536) );
  NOR2X4 U8392 ( .A(n5221), .B(n3448), .Y(n6535) );
  NOR2X4 U8393 ( .A(n5222), .B(n3448), .Y(n6538) );
  NOR2X4 U8394 ( .A(n5224), .B(n3448), .Y(n6537) );
  NOR2X4 U8395 ( .A(n5216), .B(n3460), .Y(n6544) );
  NOR2X4 U8396 ( .A(n5217), .B(n3460), .Y(n6543) );
  NOR2X4 U8397 ( .A(n5218), .B(n3460), .Y(n6546) );
  NOR2X4 U8398 ( .A(n5219), .B(n3460), .Y(n6545) );
  NOR2X4 U8399 ( .A(n5220), .B(n3460), .Y(n6548) );
  NOR2X4 U8400 ( .A(n5221), .B(n3460), .Y(n6547) );
  NOR2X4 U8401 ( .A(n5222), .B(n3460), .Y(n6550) );
  NOR2X4 U8402 ( .A(n5224), .B(n3460), .Y(n6549) );
  NOR2X4 U8403 ( .A(n5216), .B(n3459), .Y(n6556) );
  NOR2X4 U8404 ( .A(n5217), .B(n3459), .Y(n6555) );
  NOR2X4 U8405 ( .A(n5218), .B(n3459), .Y(n6558) );
  NOR2X4 U8406 ( .A(n5219), .B(n3459), .Y(n6557) );
  NOR2X4 U8407 ( .A(n5220), .B(n3459), .Y(n6560) );
  NOR2X4 U8408 ( .A(n5221), .B(n3459), .Y(n6559) );
  NOR2X4 U8409 ( .A(n5222), .B(n3459), .Y(n6562) );
  NOR2X4 U8410 ( .A(n5224), .B(n3459), .Y(n6561) );
  CMPR32X1 U8411 ( .A(n5698), .B(n4871), .C(n5256), .CO(n6117), .S(n5262) );
  ADDHXL U8412 ( .A(n6126), .B(n6127), .CO(n5256), .S(n5258) );
  OAI21XL U8413 ( .A0(n5258), .A1(n6124), .B0(n6123), .Y(n5257) );
  OAI21XL U8414 ( .A0(n5261), .A1(n5262), .B0(n5259), .Y(n5260) );
  OAI21X4 U8415 ( .A0(n5267), .A1(n6583), .B0(n5266), .Y(n6827) );
  AOI21XL U8416 ( .A0(n8259), .A1(n3395), .B0(n6827), .Y(n5271) );
  NOR2X2 U8417 ( .A(n6415), .B(n5268), .Y(n6418) );
  AOI22X4 U8418 ( .A0(N2776), .A1(n6420), .B0(n8569), .B1(n6421), .Y(n7895) );
  OAI221XL U8419 ( .A0(n7564), .A1(n5271), .B0(n8426), .B1(n8548), .C0(n5270), 
        .Y(n5272) );
  AOI22X4 U8420 ( .A0(IROM_A[5]), .A1(n5314), .B0(n5313), .B1(n8521), .Y(
        IRAM_D[7]) );
  AOI22X4 U8421 ( .A0(IROM_A[5]), .A1(n5356), .B0(n5355), .B1(n8521), .Y(
        IRAM_D[6]) );
  AOI22X4 U8422 ( .A0(IROM_A[5]), .A1(n5398), .B0(n5397), .B1(n8521), .Y(
        IRAM_D[5]) );
  AOI22X4 U8423 ( .A0(IROM_A[5]), .A1(n5440), .B0(n5439), .B1(n8521), .Y(
        IRAM_D[1]) );
  AOI22X4 U8424 ( .A0(IROM_A[5]), .A1(n5524), .B0(n5523), .B1(n8521), .Y(
        IRAM_D[0]) );
  AOI22X4 U8425 ( .A0(IROM_A[5]), .A1(n5598), .B0(n5597), .B1(n8521), .Y(
        IRAM_D[3]) );
  NAND2X2 U8426 ( .A(n8480), .B(IROM_A[4]), .Y(n6287) );
  NAND2X1 U8427 ( .A(IROM_A[5]), .B(IROM_A[3]), .Y(n7039) );
  INVX1 U8428 ( .A(n6825), .Y(n6801) );
  NOR2X4 U8429 ( .A(n6801), .B(n7029), .Y(n8295) );
  CLKINVX2 U8430 ( .A(n8295), .Y(n8329) );
  NAND2X1 U8431 ( .A(n6820), .B(n6646), .Y(n8059) );
  AOI21X1 U8432 ( .A0(n7031), .A1(n6872), .B0(n5599), .Y(n7311) );
  NOR2X1 U8433 ( .A(n7311), .B(n7306), .Y(n8333) );
  AOI21XL U8434 ( .A0(n8513), .A1(n3395), .B0(n6827), .Y(n5601) );
  CLKINVX2 U8435 ( .A(n7311), .Y(n8330) );
  OAI221XL U8436 ( .A0(n7311), .A1(n5601), .B0(n8330), .B1(n8556), .C0(n5600), 
        .Y(n5602) );
  AOI221X1 U8437 ( .A0(n6416), .A1(n5604), .B0(n6415), .B1(n5603), .C0(n6027), 
        .Y(n7973) );
  NOR2X2 U8438 ( .A(n7039), .B(n6275), .Y(n6734) );
  NOR3X2 U8439 ( .A(IROM_A[1]), .B(n8526), .C(n8519), .Y(n6779) );
  NAND2X2 U8440 ( .A(n6401), .B(n6389), .Y(n8136) );
  CLKINVX2 U8441 ( .A(n8492), .Y(n8282) );
  NAND2X2 U8442 ( .A(n8524), .B(n6742), .Y(n8125) );
  AOI21X1 U8443 ( .A0(n6734), .A1(n6779), .B0(n5606), .Y(n6273) );
  NOR2X2 U8444 ( .A(n6273), .B(n5607), .Y(n7893) );
  CMPR32X1 U8445 ( .A(DP_OP_2677J1_122_9848_n24), .B(DP_OP_2677J1_122_9848_n26), .C(n5692), .CO(n5794), .S(n5693) );
  AOI21XL U8446 ( .A0(n8492), .A1(n3375), .B0(n3437), .Y(n5702) );
  CLKINVX2 U8447 ( .A(n6273), .Y(n7890) );
  NOR2X1 U8448 ( .A(n5699), .B(n6583), .Y(n7191) );
  OAI221XL U8449 ( .A0(n6273), .A1(n5702), .B0(n7890), .B1(n8541), .C0(n5701), 
        .Y(n5703) );
  NAND2X2 U8450 ( .A(n8468), .B(n5706), .Y(n8483) );
  NAND2X1 U8451 ( .A(n8467), .B(n6984), .Y(n6668) );
  NOR2X4 U8452 ( .A(n6401), .B(n6668), .Y(n8200) );
  NOR3X2 U8453 ( .A(n8520), .B(n8526), .C(n8519), .Y(n7040) );
  AOI22X4 U8454 ( .A0(N2774), .A1(n6420), .B0(N2766), .B1(n6421), .Y(n8055) );
  CMPR32X1 U8455 ( .A(DP_OP_2677J1_122_9848_n21), .B(DP_OP_2677J1_122_9848_n23), .C(n5794), .CO(n6261), .S(n5263) );
  AOI21XL U8456 ( .A0(n8200), .A1(n7326), .B0(n3418), .Y(n5803) );
  INVX1 U8457 ( .A(n5801), .Y(n6852) );
  OAI221XL U8458 ( .A0(n5804), .A1(n5803), .B0(n8394), .B1(n8547), .C0(n5802), 
        .Y(n5805) );
  NOR3X2 U8459 ( .A(IROM_A[5]), .B(IROM_A[3]), .C(n6275), .Y(n7032) );
  NOR3X2 U8460 ( .A(IROM_A[2]), .B(n8526), .C(n8520), .Y(n7095) );
  OAI21XL U8461 ( .A0(n7029), .A1(n7033), .B0(n8446), .Y(n5811) );
  NAND2X2 U8462 ( .A(n6699), .B(n5929), .Y(n8406) );
  AOI21X1 U8463 ( .A0(n7032), .A1(n7095), .B0(n5810), .Y(n8034) );
  NOR2X2 U8464 ( .A(n8034), .B(n5811), .Y(n8451) );
  AOI22X1 U8465 ( .A0(N2772), .A1(n6420), .B0(n8567), .B1(n6421), .Y(n5812) );
  AOI21XL U8466 ( .A0(n8032), .A1(n3350), .B0(n3440), .Y(n5905) );
  CLKINVX2 U8467 ( .A(n8034), .Y(n8448) );
  AOI22X4 U8468 ( .A0(N2772), .A1(n6421), .B0(n8567), .B1(n6420), .Y(n7740) );
  OAI221XL U8469 ( .A0(n8034), .A1(n5905), .B0(n8448), .B1(n8551), .C0(n5904), 
        .Y(n5906) );
  NAND2X2 U8470 ( .A(n6030), .B(n3453), .Y(n8159) );
  NOR2X1 U8471 ( .A(n6902), .B(n6800), .Y(n6791) );
  NAND2X1 U8472 ( .A(n8524), .B(n6791), .Y(n7864) );
  CLKINVX2 U8473 ( .A(n7935), .Y(n8160) );
  AOI21XL U8474 ( .A0(n8228), .A1(n3395), .B0(n6827), .Y(n5912) );
  OAI221XL U8475 ( .A0(n7935), .A1(n5912), .B0(n8160), .B1(n8542), .C0(n5911), 
        .Y(n5913) );
  INVX1 U8476 ( .A(n3455), .Y(n8023) );
  NOR2X2 U8477 ( .A(n5914), .B(n8483), .Y(n7513) );
  NOR2X2 U8478 ( .A(n5919), .B(n5916), .Y(n7701) );
  AOI21XL U8479 ( .A0(n3455), .A1(n6880), .B0(n6827), .Y(n5918) );
  OAI221XL U8480 ( .A0(n5919), .A1(n5918), .B0(n7698), .B1(n8539), .C0(n5917), 
        .Y(n5920) );
  NOR2X1 U8481 ( .A(n6800), .B(n6776), .Y(n6721) );
  NAND2X2 U8482 ( .A(n8524), .B(n3413), .Y(n7907) );
  AOI21XL U8483 ( .A0(n6401), .A1(n6625), .B0(n8501), .Y(n5923) );
  NOR3X2 U8484 ( .A(IROM_A[5]), .B(n6287), .C(n8522), .Y(n6760) );
  NOR2X4 U8485 ( .A(n6401), .B(n6634), .Y(n8499) );
  AOI21X1 U8486 ( .A0(n6760), .A1(n7095), .B0(n5922), .Y(n6980) );
  CLKINVX2 U8487 ( .A(n6980), .Y(n8178) );
  AOI21XL U8488 ( .A0(n8501), .A1(n3375), .B0(n3437), .Y(n5926) );
  NAND2X1 U8489 ( .A(op4[3]), .B(n6721), .Y(n8177) );
  OAI221XL U8490 ( .A0(n6980), .A1(n5926), .B0(n8178), .B1(n8562), .C0(n5925), 
        .Y(n5927) );
  NOR3X2 U8491 ( .A(IROM_A[1]), .B(IROM_A[2]), .C(n8526), .Y(n6871) );
  OAI221X4 U8492 ( .A0(n6416), .A1(N2757), .B0(n6415), .B1(N2781), .C0(n6414), 
        .Y(n7307) );
  AOI21XL U8493 ( .A0(n3361), .A1(n6970), .B0(n3464), .Y(n6022) );
  AOI22X4 U8494 ( .A0(N2773), .A1(n6421), .B0(N2765), .B1(n6420), .Y(n7963) );
  AOI22X4 U8495 ( .A0(N2773), .A1(n6420), .B0(N2765), .B1(n6421), .Y(n7956) );
  AOI21XL U8496 ( .A0(n8301), .A1(n7326), .B0(n3418), .Y(n6025) );
  OAI221XL U8497 ( .A0(n6980), .A1(n6025), .B0(n8178), .B1(n8561), .C0(n6024), 
        .Y(n6026) );
  NOR2X1 U8498 ( .A(n6747), .B(n7034), .Y(n6786) );
  NAND2X1 U8499 ( .A(op4[3]), .B(n6786), .Y(n7925) );
  AOI21X1 U8500 ( .A0(n7031), .A1(n6734), .B0(n6031), .Y(n6884) );
  CMPR32X1 U8501 ( .A(DP_OP_2677J1_122_9848_n27), .B(n6117), .C(n6116), .CO(
        n5692), .S(n6118) );
  AOI21XL U8502 ( .A0(n5908), .A1(n3356), .B0(n3439), .Y(n6129) );
  CLKINVX2 U8503 ( .A(n6884), .Y(n8269) );
  NOR2X1 U8504 ( .A(n6125), .B(n6583), .Y(n6145) );
  OAI221XL U8505 ( .A0(n6884), .A1(n6129), .B0(n8269), .B1(n8544), .C0(n6128), 
        .Y(n6130) );
  NOR2X4 U8506 ( .A(n6131), .B(n6650), .Y(n8343) );
  NAND2X2 U8507 ( .A(n8467), .B(n6825), .Y(n8076) );
  NOR3X2 U8508 ( .A(IROM_A[1]), .B(IROM_A[0]), .C(IROM_A[2]), .Y(n6688) );
  AOI21X1 U8509 ( .A0(n6688), .A1(n6872), .B0(n6132), .Y(n8079) );
  AOI21XL U8510 ( .A0(n8343), .A1(n7326), .B0(n3418), .Y(n6134) );
  AOI21XL U8511 ( .A0(n6401), .A1(n6720), .B0(n8499), .Y(n7972) );
  NOR3X2 U8512 ( .A(IROM_A[1]), .B(IROM_A[0]), .C(n8519), .Y(n7008) );
  CLKINVX3 U8513 ( .A(n7826), .Y(n8289) );
  CLKINVX2 U8514 ( .A(n7978), .Y(n8154) );
  AOI21XL U8515 ( .A0(n8499), .A1(n3360), .B0(n3439), .Y(n6140) );
  OAI221XL U8516 ( .A0(n7978), .A1(n6140), .B0(n8154), .B1(n8560), .C0(n6139), 
        .Y(n6141) );
  INVX1 U8517 ( .A(n3449), .Y(n6748) );
  AOI21XL U8518 ( .A0(n6401), .A1(n6338), .B0(n7898), .Y(n7983) );
  CLKINVX2 U8519 ( .A(n7987), .Y(n8143) );
  NAND2X1 U8520 ( .A(n3449), .B(n6984), .Y(n6665) );
  AOI21XL U8521 ( .A0(n8114), .A1(n8141), .B0(n3439), .Y(n6148) );
  OAI221XL U8522 ( .A0(n7987), .A1(n6148), .B0(n8143), .B1(n8564), .C0(n6147), 
        .Y(n6149) );
  NOR2X4 U8523 ( .A(n6401), .B(n6650), .Y(n8215) );
  NOR3X2 U8524 ( .A(IROM_A[3]), .B(n8521), .C(n6287), .Y(n6904) );
  AOI21XL U8525 ( .A0(n8215), .A1(n3356), .B0(n3439), .Y(n6153) );
  OAI221XL U8526 ( .A0(n6154), .A1(n6153), .B0(n8240), .B1(n8559), .C0(n6152), 
        .Y(n6155) );
  AOI21XL U8527 ( .A0(n8214), .A1(n7581), .B0(n3440), .Y(n6157) );
  OAI221XL U8528 ( .A0(n6884), .A1(n6157), .B0(n8269), .B1(n8543), .C0(n6156), 
        .Y(n6158) );
  AOI21XL U8529 ( .A0(n3353), .A1(n3383), .B0(n3440), .Y(n6162) );
  OAI221XL U8530 ( .A0(n6163), .A1(n6162), .B0(n8172), .B1(n8563), .C0(n6161), 
        .Y(n6164) );
  AOI21XL U8531 ( .A0(n3353), .A1(n3380), .B0(n3440), .Y(n6169) );
  OAI221XL U8532 ( .A0(n6170), .A1(n6169), .B0(n8166), .B1(n8545), .C0(n6168), 
        .Y(n6171) );
  OAI21XL U8533 ( .A0(N2783), .A1(n6417), .B0(n6414), .Y(n6172) );
  NOR2X4 U8534 ( .A(n6748), .B(n6766), .Y(n8260) );
  NOR2X2 U8535 ( .A(n6269), .B(n6175), .Y(n8094) );
  OAI21X4 U8536 ( .A0(n6266), .A1(n6583), .B0(n6265), .Y(n6403) );
  AOI21XL U8537 ( .A0(n3389), .A1(n8417), .B0(n6403), .Y(n6268) );
  AOI22X4 U8538 ( .A0(N2775), .A1(n6420), .B0(n8568), .B1(n6421), .Y(n8447) );
  AOI22X1 U8539 ( .A0(N2775), .A1(n6421), .B0(n8568), .B1(n6420), .Y(n8268) );
  OAI221XL U8540 ( .A0(n6269), .A1(n6268), .B0(n8091), .B1(n8549), .C0(n6267), 
        .Y(n6270) );
  AOI21XL U8541 ( .A0(n3389), .A1(n7888), .B0(n6403), .Y(n6272) );
  OAI221XL U8542 ( .A0(n6273), .A1(n6272), .B0(n7890), .B1(n8540), .C0(n6271), 
        .Y(n6274) );
  NOR3X2 U8543 ( .A(IROM_A[3]), .B(n8521), .C(n6275), .Y(n6994) );
  AOI21X1 U8544 ( .A0(n6994), .A1(n7095), .B0(n6276), .Y(n6279) );
  NOR3X2 U8545 ( .A(n3413), .B(n8499), .C(n6279), .Y(n7910) );
  AOI21XL U8546 ( .A0(n3389), .A1(n8501), .B0(n6403), .Y(n6278) );
  OAI221XL U8547 ( .A0(n6279), .A1(n6278), .B0(n8507), .B1(n8546), .C0(n6277), 
        .Y(n6280) );
  AOI21XL U8548 ( .A0(n8295), .A1(n3395), .B0(n6827), .Y(n6284) );
  OAI221XL U8549 ( .A0(n6285), .A1(n6284), .B0(n7349), .B1(n8558), .C0(n6283), 
        .Y(n6286) );
  NOR3X2 U8550 ( .A(IROM_A[5]), .B(IROM_A[3]), .C(n6287), .Y(n6986) );
  AOI21X1 U8551 ( .A0(n6986), .A1(n3410), .B0(n6288), .Y(n6294) );
  AOI211X2 U8552 ( .A0(n6984), .A1(n3400), .B0(n3382), .C0(n6294), .Y(n7922)
         );
  AOI21XL U8553 ( .A0(n8287), .A1(n3349), .B0(n6403), .Y(n6293) );
  OAI221XL U8554 ( .A0(n6294), .A1(n6293), .B0(n7919), .B1(n8565), .C0(n6292), 
        .Y(n6295) );
  INVXL U8555 ( .A(n6386), .Y(n6318) );
  OAI21XL U8556 ( .A0(n7033), .A1(n6318), .B0(n6902), .Y(n6302) );
  NOR2X1 U8557 ( .A(cmd_reg[2]), .B(n6304), .Y(n6301) );
  OAI21XL U8558 ( .A0(n6710), .A1(n6299), .B0(n6747), .Y(n6300) );
  AOI22XL U8559 ( .A0(n6303), .A1(n6302), .B0(n6301), .B1(n6300), .Y(n6306) );
  OR3XL U8560 ( .A(n6304), .B(cmd_reg[2]), .C(n6312), .Y(n6319) );
  INVXL U8561 ( .A(n6385), .Y(n6305) );
  CLKINVX3 U8562 ( .A(reset), .Y(n8588) );
  CLKINVX3 U8563 ( .A(reset), .Y(n8589) );
  CLKINVX3 U8564 ( .A(reset), .Y(n8590) );
  CLKINVX3 U8565 ( .A(reset), .Y(n8591) );
  CLKINVX3 U8566 ( .A(reset), .Y(n8592) );
  CLKINVX3 U8567 ( .A(reset), .Y(n8593) );
  CLKINVX3 U8568 ( .A(reset), .Y(n8582) );
  CLKINVX3 U8569 ( .A(reset), .Y(n8584) );
  CLKINVX3 U8570 ( .A(reset), .Y(n8581) );
  CLKINVX3 U8571 ( .A(reset), .Y(n8585) );
  CLKINVX3 U8572 ( .A(reset), .Y(n8586) );
  CLKINVX3 U8573 ( .A(reset), .Y(n8580) );
  CLKINVX3 U8574 ( .A(reset), .Y(n8587) );
  CLKINVX3 U8575 ( .A(reset), .Y(n8597) );
  CLKINVX3 U8576 ( .A(reset), .Y(n8601) );
  CLKINVX3 U8577 ( .A(reset), .Y(n8598) );
  CLKINVX3 U8578 ( .A(reset), .Y(n8573) );
  CLKINVX3 U8579 ( .A(reset), .Y(n8600) );
  CLKINVX3 U8580 ( .A(reset), .Y(n8572) );
  CLKINVX3 U8581 ( .A(reset), .Y(n8599) );
  CLKINVX3 U8582 ( .A(reset), .Y(n8594) );
  CLKINVX3 U8583 ( .A(reset), .Y(n8575) );
  CLKINVX3 U8584 ( .A(reset), .Y(n8602) );
  CLKINVX3 U8585 ( .A(reset), .Y(n8570) );
  CLKINVX3 U8586 ( .A(reset), .Y(n8596) );
  CLKINVX3 U8587 ( .A(reset), .Y(n8574) );
  INVXL U8588 ( .A(n8466), .Y(n8472) );
  NOR2X1 U8589 ( .A(n8532), .B(n6311), .Y(n8473) );
  NAND2XL U8590 ( .A(n8473), .B(n8529), .Y(n8469) );
  AOI21XL U8591 ( .A0(n8472), .A1(n8469), .B0(n6312), .Y(n6315) );
  NAND2XL U8592 ( .A(op2[0]), .B(n6748), .Y(n8471) );
  OAI21XL U8593 ( .A0(n8473), .A1(n8466), .B0(n6313), .Y(n8475) );
  INVXL U8594 ( .A(n8475), .Y(n8470) );
  OAI22XL U8595 ( .A0(n8470), .A1(n8529), .B0(n8483), .B1(n8482), .Y(n6314) );
  AOI21XL U8596 ( .A0(n6315), .A1(n8471), .B0(n6314), .Y(n3324) );
  INVXL U8597 ( .A(n6316), .Y(n6321) );
  AOI31XL U8598 ( .A0(cs[0]), .A1(cmd_valid), .A2(n8533), .B0(n6322), .Y(n3327) );
  INVXL U8599 ( .A(n8489), .Y(n8460) );
  AOI21XL U8600 ( .A0(n3361), .A1(n6592), .B0(n3464), .Y(n6326) );
  CLKINVX2 U8601 ( .A(n8141), .Y(n8275) );
  CLKINVX2 U8602 ( .A(n8259), .Y(n8425) );
  NAND2XL U8603 ( .A(n6665), .B(n8425), .Y(n6682) );
  AOI22X1 U8604 ( .A0(n6986), .A1(n6871), .B0(n3398), .B1(n6338), .Y(n6683) );
  NAND2XL U8605 ( .A(n8351), .B(n6758), .Y(n6677) );
  CLKINVX3 U8606 ( .A(n7513), .Y(n8381) );
  NAND3XL U8607 ( .A(n8023), .B(n8381), .C(n8165), .Y(n6672) );
  NOR2X2 U8608 ( .A(n6802), .B(n3438), .Y(n8038) );
  AOI21XL U8609 ( .A0(n6353), .A1(n6780), .B0(n8038), .Y(n6975) );
  CLKINVX3 U8610 ( .A(n8038), .Y(n8432) );
  NOR2X4 U8611 ( .A(n6777), .B(n6767), .Y(n8385) );
  AOI21XL U8612 ( .A0(n3369), .A1(n6975), .B0(n6403), .Y(n6363) );
  OAI221XL U8613 ( .A0(n6978), .A1(n6363), .B0(n8086), .B1(n8550), .C0(n6362), 
        .Y(n6364) );
  AOI21XL U8614 ( .A0(n8519), .A1(n8464), .B0(n8487), .Y(n6381) );
  OAI21XL U8615 ( .A0(n7033), .A1(n6384), .B0(n6383), .Y(n6387) );
  NOR2X1 U8616 ( .A(n3423), .B(n6950), .Y(n7486) );
  AOI21XL U8617 ( .A0(n8315), .A1(n7326), .B0(n3418), .Y(n6392) );
  CLKINVX2 U8618 ( .A(n3423), .Y(n7483) );
  AOI21XL U8619 ( .A0(n7888), .A1(n3395), .B0(n6827), .Y(n6395) );
  AOI21XL U8620 ( .A0(n6401), .A1(n6398), .B0(n3376), .Y(n6400) );
  CLKINVX2 U8621 ( .A(n3425), .Y(n6957) );
  NAND2X2 U8622 ( .A(n6401), .B(n6742), .Y(n8070) );
  OAI21XL U8623 ( .A0(n8447), .A1(n8070), .B0(n6402), .Y(n6405) );
  OAI21XL U8624 ( .A0(n8372), .A1(n7002), .B0(n3347), .Y(n6410) );
  OAI21XL U8625 ( .A0(n6407), .A1(n8406), .B0(n6408), .Y(n6409) );
  OAI21XL U8626 ( .A0(n8199), .A1(n6950), .B0(n3347), .Y(n6413) );
  OAI21XL U8627 ( .A0(n6407), .A1(n8289), .B0(n6411), .Y(n6412) );
  OAI221X4 U8628 ( .A0(n6416), .A1(N2755), .B0(n6415), .B1(N2779), .C0(n6414), 
        .Y(n7578) );
  AOI22X4 U8629 ( .A0(N2771), .A1(n6420), .B0(n3442), .B1(n6421), .Y(n7570) );
  INVX1 U8630 ( .A(n8362), .Y(n8153) );
  NOR2X2 U8631 ( .A(n6419), .B(n6583), .Y(n6973) );
  AOI22X1 U8632 ( .A0(N2771), .A1(n6421), .B0(n3442), .B1(n6420), .Y(n6893) );
  OAI21XL U8633 ( .A0(n7570), .A1(n8153), .B0(n6422), .Y(n6588) );
  CMPR32X1 U8634 ( .A(DP_OP_2677J1_122_9848_n11), .B(DP_OP_2677J1_122_9848_n10), .C(n6575), .CO(n6576), .S(n5898) );
  OAI221XL U8635 ( .A0(in_valid), .A1(IRAM_D[7]), .B0(n8523), .B1(IROM_Q[7]), 
        .C0(n8480), .Y(n6582) );
  OAI21XL U8636 ( .A0(n3394), .A1(n8351), .B0(n6589), .Y(n6591) );
  OAI21XL U8637 ( .A0(n7570), .A1(n8136), .B0(n6593), .Y(n6595) );
  OAI21XL U8638 ( .A0(n3394), .A1(n7907), .B0(n6596), .Y(n6598) );
  OAI21XL U8639 ( .A0(n3394), .A1(n8165), .B0(n6599), .Y(n6601) );
  OAI21XL U8640 ( .A0(n3394), .A1(n8171), .B0(n6602), .Y(n6604) );
  OAI21XL U8641 ( .A0(n3394), .A1(n8329), .B0(n6605), .Y(n6607) );
  OAI21XL U8642 ( .A0(n3394), .A1(n8159), .B0(n6608), .Y(n6610) );
  OAI21XL U8643 ( .A0(n7570), .A1(n8393), .B0(n6611), .Y(n6613) );
  OAI21XL U8644 ( .A0(n7570), .A1(n8209), .B0(n6617), .Y(n6619) );
  OAI21XL U8645 ( .A0(n3394), .A1(n8184), .B0(n6622), .Y(n6624) );
  OAI21XL U8646 ( .A0(n7570), .A1(n8304), .B0(n6628), .Y(n6630) );
  OAI21XL U8647 ( .A0(n7570), .A1(n8289), .B0(n6635), .Y(n6637) );
  NAND2XL U8648 ( .A(n7918), .B(n3397), .Y(n6640) );
  OAI21XL U8649 ( .A0(n7570), .A1(n3397), .B0(n6642), .Y(n6645) );
  OAI21XL U8650 ( .A0(n3393), .A1(n8310), .B0(n6652), .Y(n6654) );
  OAI21XL U8651 ( .A0(n3394), .A1(n3405), .B0(n6659), .Y(n6661) );
  OAI21XL U8652 ( .A0(n6893), .A1(n8076), .B0(n6662), .Y(n6664) );
  OAI21XL U8653 ( .A0(n3393), .A1(n8393), .B0(n6669), .Y(n6671) );
  OAI21XL U8654 ( .A0(n6893), .A1(n8381), .B0(n6674), .Y(n6676) );
  OAI21XL U8655 ( .A0(n7570), .A1(n8351), .B0(n6679), .Y(n6681) );
  OAI21XL U8656 ( .A0(n3393), .A1(n7684), .B0(n6684), .Y(n6686) );
  NOR2X2 U8657 ( .A(n6691), .B(n6689), .Y(n8279) );
  OAI21XL U8658 ( .A0(n7570), .A1(n8275), .B0(n6690), .Y(n6693) );
  OAI21XL U8659 ( .A0(n3394), .A1(n8267), .B0(n6694), .Y(n6696) );
  AOI22X1 U8660 ( .A0(n6904), .A1(n7008), .B0(n3398), .B1(n6698), .Y(n6701) );
  NOR3X2 U8661 ( .A(n6791), .B(n8492), .C(n6701), .Y(n8286) );
  NAND2X1 U8662 ( .A(n6825), .B(n6699), .Y(n7455) );
  OAI21XL U8663 ( .A0(n3394), .A1(n7455), .B0(n6700), .Y(n6703) );
  AOI22X1 U8664 ( .A0(n6779), .A1(n7096), .B0(n3398), .B1(n6704), .Y(n6707) );
  CLKINVX3 U8665 ( .A(n8302), .Y(n8387) );
  NOR2X2 U8666 ( .A(n6707), .B(n6705), .Y(n8391) );
  OAI21XL U8667 ( .A0(n3394), .A1(n8387), .B0(n6706), .Y(n6709) );
  AOI22X1 U8668 ( .A0(n6779), .A1(n6760), .B0(n3398), .B1(n6711), .Y(n6714) );
  NOR2X2 U8669 ( .A(n6714), .B(n6712), .Y(n8293) );
  OAI21XL U8670 ( .A0(n3394), .A1(n8289), .B0(n6713), .Y(n6716) );
  OAI21XL U8671 ( .A0(n3394), .A1(n8125), .B0(n6717), .Y(n6719) );
  OAI21XL U8672 ( .A0(n7570), .A1(n8387), .B0(n6722), .Y(n6725) );
  NOR2X4 U8673 ( .A(n6728), .B(n8483), .Y(n8356) );
  CLKINVX2 U8674 ( .A(n8356), .Y(n8130) );
  NOR2X2 U8675 ( .A(n3412), .B(n6729), .Y(n8321) );
  OAI21XL U8676 ( .A0(n7570), .A1(n8130), .B0(n6730), .Y(n6732) );
  AOI21X1 U8677 ( .A0(n6871), .A1(n6734), .B0(n6733), .Y(n7940) );
  NOR2X2 U8678 ( .A(n7940), .B(n6735), .Y(n8314) );
  OAI21XL U8679 ( .A0(n3394), .A1(n8310), .B0(n6736), .Y(n6738) );
  OAI21XL U8680 ( .A0(n3394), .A1(n8282), .B0(n6739), .Y(n6741) );
  AOI22X1 U8681 ( .A0(n6904), .A1(n3410), .B0(n3398), .B1(n6819), .Y(n6744) );
  NOR3X2 U8682 ( .A(n6742), .B(n7513), .C(n6744), .Y(n8339) );
  OAI21XL U8683 ( .A0(n7570), .A1(n8381), .B0(n6743), .Y(n6746) );
  AOI211X2 U8684 ( .A0(n3449), .A1(n6991), .B0(n6143), .C0(n6752), .Y(n8355)
         );
  OAI21XL U8685 ( .A0(n3394), .A1(n8349), .B0(n6751), .Y(n6754) );
  OAI21XL U8686 ( .A0(n7570), .A1(n7975), .B0(n6755), .Y(n6757) );
  NAND2XL U8687 ( .A(n8130), .B(n3397), .Y(n6761) );
  OAI21XL U8688 ( .A0(n3393), .A1(n3397), .B0(n6762), .Y(n6765) );
  OAI21XL U8689 ( .A0(n3393), .A1(n8454), .B0(n6769), .Y(n6772) );
  OAI21XL U8690 ( .A0(n3394), .A1(n7918), .B0(n6773), .Y(n6775) );
  AOI211X2 U8691 ( .A0(n6984), .A1(n6780), .B0(n3384), .C0(n6782), .Y(n8367)
         );
  OAI21XL U8692 ( .A0(n3393), .A1(n8387), .B0(n6781), .Y(n6784) );
  NOR3X2 U8693 ( .A(n6786), .B(n8501), .C(n6785), .Y(n7929) );
  OAI21XL U8694 ( .A0(n7570), .A1(n7907), .B0(n6788), .Y(n6790) );
  OAI21XL U8695 ( .A0(n6792), .A1(n6791), .B0(op4[3]), .Y(n6795) );
  OAI21XL U8696 ( .A0(n7740), .A1(n8446), .B0(n6796), .Y(n6799) );
  AOI22X1 U8697 ( .A0(n6872), .A1(n7095), .B0(n3398), .B1(n6803), .Y(n6806) );
  CLKINVX3 U8698 ( .A(n8511), .Y(n8412) );
  NOR2X2 U8699 ( .A(n6806), .B(n6804), .Y(n8300) );
  OAI21XL U8700 ( .A0(n7740), .A1(n8412), .B0(n6805), .Y(n6808) );
  OAI21XL U8701 ( .A0(n3419), .A1(n8446), .B0(n6809), .Y(n6812) );
  OAI21XL U8702 ( .A0(n3385), .A1(n8329), .B0(n6813), .Y(n6815) );
  OAI21XL U8703 ( .A0(n3419), .A1(n8412), .B0(n6816), .Y(n6818) );
  NAND2X1 U8704 ( .A(n6825), .B(n6992), .Y(n8440) );
  OAI21XL U8705 ( .A0(n3372), .A1(n8432), .B0(n6826), .Y(n6829) );
  OAI21XL U8706 ( .A0(n7895), .A1(n8070), .B0(n6830), .Y(n6832) );
  OAI21XL U8707 ( .A0(n3372), .A1(n8412), .B0(n6833), .Y(n6835) );
  OAI21XL U8708 ( .A0(n7963), .A1(n8446), .B0(n6836), .Y(n6839) );
  OAI21XL U8709 ( .A0(n7963), .A1(n8432), .B0(n6840), .Y(n6842) );
  OAI21XL U8710 ( .A0(n7956), .A1(n8070), .B0(n6843), .Y(n6845) );
  OAI21XL U8711 ( .A0(n7963), .A1(n8412), .B0(n6846), .Y(n6848) );
  OAI21XL U8712 ( .A0(n7963), .A1(n8070), .B0(n6849), .Y(n6851) );
  OAI21XL U8713 ( .A0(n3370), .A1(n8432), .B0(n6853), .Y(n6857) );
  OAI21XL U8714 ( .A0(n3370), .A1(n8446), .B0(n6858), .Y(n6860) );
  OAI21XL U8715 ( .A0(n8055), .A1(n8070), .B0(n6861), .Y(n6863) );
  OAI21XL U8716 ( .A0(n8055), .A1(n8329), .B0(n6864), .Y(n6866) );
  OAI21XL U8717 ( .A0(n3370), .A1(n8412), .B0(n6867), .Y(n6869) );
  INVX1 U8718 ( .A(n8343), .Y(n8217) );
  AOI22X1 U8719 ( .A0(n6872), .A1(n6871), .B0(n3398), .B1(n6870), .Y(n6875) );
  NAND2XL U8720 ( .A(n3405), .B(n8217), .Y(n6873) );
  NOR3X2 U8721 ( .A(n8182), .B(n6875), .C(n6873), .Y(n8348) );
  OAI21XL U8722 ( .A0(n3370), .A1(n8370), .B0(n6874), .Y(n6877) );
  OAI21XL U8723 ( .A0(n7773), .A1(n7925), .B0(n6881), .Y(n6882) );
  OAI21XL U8724 ( .A0(n7570), .A1(n8070), .B0(n6888), .Y(n6890) );
  OAI21XL U8725 ( .A0(n6893), .A1(n8446), .B0(n6892), .Y(n6895) );
  OAI21XL U8726 ( .A0(n3394), .A1(n8432), .B0(n6896), .Y(n6898) );
  OAI21XL U8727 ( .A0(n3394), .A1(n8412), .B0(n6899), .Y(n6901) );
  OAI21XL U8728 ( .A0(n8483), .A1(n6902), .B0(n8076), .Y(n6905) );
  NOR2X2 U8729 ( .A(n8380), .B(n6905), .Y(n8384) );
  OAI21XL U8730 ( .A0(n3393), .A1(n8381), .B0(n6906), .Y(n6908) );
  OAI21XL U8731 ( .A0(n3394), .A1(n8323), .B0(n6909), .Y(n6911) );
  OAI21XL U8732 ( .A0(n7570), .A1(n8329), .B0(n6912), .Y(n6914) );
  OAI21XL U8733 ( .A0(n6893), .A1(n8370), .B0(n6915), .Y(n6917) );
  OAI21XL U8734 ( .A0(n3359), .A1(n8446), .B0(n6918), .Y(n6921) );
  OAI21XL U8735 ( .A0(n3359), .A1(n8432), .B0(n6922), .Y(n6924) );
  OAI21XL U8736 ( .A0(n3374), .A1(n8381), .B0(n6925), .Y(n6927) );
  OAI21XL U8737 ( .A0(n3359), .A1(n8323), .B0(n6928), .Y(n6930) );
  OAI21XL U8738 ( .A0(n3421), .A1(n8329), .B0(n6931), .Y(n6933) );
  OAI21XL U8739 ( .A0(n3359), .A1(n8412), .B0(n6937), .Y(n6939) );
  OAI21XL U8740 ( .A0(n3359), .A1(n8070), .B0(n6940), .Y(n6942) );
  OAI21XL U8741 ( .A0(n3359), .A1(n8370), .B0(n6944), .Y(n6946) );
  OAI21XL U8742 ( .A0(n8509), .A1(n6950), .B0(n3365), .Y(n6954) );
  OAI21XL U8743 ( .A0(n3392), .A1(n8289), .B0(n6952), .Y(n6953) );
  OAI21XL U8744 ( .A0(n3396), .A1(n8070), .B0(n3365), .Y(n6958) );
  OAI21XL U8745 ( .A0(n8069), .A1(n8509), .B0(n6955), .Y(n6956) );
  OAI21XL U8746 ( .A0(n3385), .A1(n8202), .B0(n3367), .Y(n6990) );
  OAI21XL U8747 ( .A0(n3390), .A1(n7566), .B0(n6988), .Y(n6989) );
  AOI21X1 U8748 ( .A0(n7040), .A1(n6994), .B0(n6993), .Y(n8026) );
  OAI21XL U8749 ( .A0(n3419), .A1(n8023), .B0(n3367), .Y(n6997) );
  CLKINVX2 U8750 ( .A(n8026), .Y(n8131) );
  OAI21XL U8751 ( .A0(n3390), .A1(n7577), .B0(n6995), .Y(n6996) );
  OAI21XL U8752 ( .A0(n3390), .A1(n6998), .B0(n3367), .Y(n7001) );
  OAI21XL U8753 ( .A0(n8111), .A1(n3399), .B0(n6999), .Y(n7000) );
  OAI21XL U8754 ( .A0(n7570), .A1(n7995), .B0(n7004), .Y(n7006) );
  OAI21XL U8755 ( .A0(n3393), .A1(n8446), .B0(n7011), .Y(n7013) );
  AOI21X1 U8756 ( .A0(n7032), .A1(n3410), .B0(n7015), .Y(n7747) );
  NOR3X2 U8757 ( .A(n8430), .B(n7747), .C(n7016), .Y(n8436) );
  OAI21XL U8758 ( .A0(n8432), .A1(n3393), .B0(n7017), .Y(n7019) );
  NAND2XL U8759 ( .A(n8419), .B(n8184), .Y(n7021) );
  OAI21XL U8760 ( .A0(n3393), .A1(n8419), .B0(n7022), .Y(n7025) );
  OAI21XL U8761 ( .A0(n3394), .A1(n8393), .B0(n7026), .Y(n7028) );
  OAI21XL U8762 ( .A0(n7034), .A1(n7033), .B0(n8412), .Y(n8508) );
  OAI21XL U8763 ( .A0(n3394), .A1(n8101), .B0(n7036), .Y(n7038) );
  NAND2XL U8764 ( .A(n8419), .B(n8440), .Y(n7044) );
  OAI21XL U8765 ( .A0(n7570), .A1(n8323), .B0(n7045), .Y(n7048) );
  OAI21XL U8766 ( .A0(n3393), .A1(n8412), .B0(n7049), .Y(n7051) );
  OAI21XL U8767 ( .A0(n3394), .A1(n7684), .B0(n7052), .Y(n7054) );
  OAI21XL U8768 ( .A0(n3374), .A1(n8130), .B0(n7062), .Y(n7064) );
  OAI21XL U8769 ( .A0(n3391), .A1(n8130), .B0(n7065), .Y(n7067) );
  OAI21XL U8770 ( .A0(n3421), .A1(n8136), .B0(n7069), .Y(n7071) );
  INVX1 U8771 ( .A(n7566), .Y(n8151) );
  OAI21XL U8772 ( .A0(n3359), .A1(n3397), .B0(n7072), .Y(n7074) );
  OAI21XL U8773 ( .A0(n7956), .A1(n8153), .B0(n7075), .Y(n7077) );
  OAI21XL U8774 ( .A0(n7963), .A1(n3397), .B0(n7079), .Y(n7081) );
  OAI21XL U8775 ( .A0(n7963), .A1(n8351), .B0(n7082), .Y(n7084) );
  OAI21XL U8776 ( .A0(n7956), .A1(n7864), .B0(n7085), .Y(n7087) );
  OAI21XL U8777 ( .A0(n7963), .A1(n8165), .B0(n7088), .Y(n7090) );
  OAI21XL U8778 ( .A0(n3359), .A1(n8165), .B0(n7091), .Y(n7093) );
  OAI21XL U8779 ( .A0(n3421), .A1(n8406), .B0(n7098), .Y(n7100) );
  OAI21XL U8780 ( .A0(n7956), .A1(n8406), .B0(n7101), .Y(n7103) );
  OAI21XL U8781 ( .A0(n7956), .A1(n8393), .B0(n7104), .Y(n7106) );
  OAI21XL U8782 ( .A0(n3359), .A1(n8159), .B0(n7107), .Y(n7109) );
  OAI21XL U8783 ( .A0(n3359), .A1(n8171), .B0(n7110), .Y(n7112) );
  OAI21XL U8784 ( .A0(n3421), .A1(n8393), .B0(n7113), .Y(n7115) );
  OAI21XL U8785 ( .A0(n7963), .A1(n8171), .B0(n7116), .Y(n7118) );
  OAI21XL U8786 ( .A0(n3421), .A1(n8370), .B0(n7119), .Y(n7121) );
  OAI21XL U8787 ( .A0(n3391), .A1(n8209), .B0(n7122), .Y(n7124) );
  OAI21XL U8788 ( .A0(n7963), .A1(n8217), .B0(n7125), .Y(n7127) );
  OAI21XL U8789 ( .A0(n7956), .A1(n8209), .B0(n7128), .Y(n7130) );
  OAI21XL U8790 ( .A0(n3421), .A1(n8209), .B0(n7131), .Y(n7133) );
  OAI21XL U8791 ( .A0(n7963), .A1(n8184), .B0(n7134), .Y(n7136) );
  OAI21XL U8792 ( .A0(n7956), .A1(n7684), .B0(n7137), .Y(n7139) );
  OAI21XL U8793 ( .A0(n3421), .A1(n8289), .B0(n7140), .Y(n7142) );
  OAI21XL U8794 ( .A0(n3421), .A1(n7684), .B0(n7143), .Y(n7145) );
  OAI21XL U8795 ( .A0(n3421), .A1(n8304), .B0(n7146), .Y(n7148) );
  OAI21XL U8796 ( .A0(n7956), .A1(n3397), .B0(n7149), .Y(n7151) );
  OAI21XL U8797 ( .A0(n7956), .A1(n8159), .B0(n7152), .Y(n7154) );
  OAI21XL U8798 ( .A0(n3391), .A1(n7975), .B0(n7155), .Y(n7157) );
  OAI21XL U8799 ( .A0(n3391), .A1(n8165), .B0(n7158), .Y(n7160) );
  OAI21XL U8800 ( .A0(n3359), .A1(n8217), .B0(n7161), .Y(n7163) );
  OAI21XL U8801 ( .A0(n7963), .A1(n8381), .B0(n7164), .Y(n7166) );
  OAI21XL U8802 ( .A0(n3421), .A1(n3397), .B0(n7167), .Y(n7169) );
  OAI21XL U8803 ( .A0(n3359), .A1(n8076), .B0(n7170), .Y(n7172) );
  OAI21XL U8804 ( .A0(n3359), .A1(n8381), .B0(n7173), .Y(n7175) );
  OAI21XL U8805 ( .A0(n3359), .A1(n3405), .B0(n7176), .Y(n7178) );
  OAI21XL U8806 ( .A0(n3421), .A1(n8351), .B0(n7179), .Y(n7181) );
  OAI21XL U8807 ( .A0(n3421), .A1(n8425), .B0(n7182), .Y(n7184) );
  OAI21XL U8808 ( .A0(n7956), .A1(n7995), .B0(n7185), .Y(n7187) );
  OAI21XL U8809 ( .A0(n3421), .A1(n7995), .B0(n7188), .Y(n7190) );
  OAI21XL U8810 ( .A0(n3374), .A1(n7864), .B0(n7192), .Y(n7194) );
  OAI21XL U8811 ( .A0(n7963), .A1(n8267), .B0(n7195), .Y(n7197) );
  OAI21XL U8812 ( .A0(n3359), .A1(n8267), .B0(n7198), .Y(n7200) );
  OAI21XL U8813 ( .A0(n7956), .A1(n8275), .B0(n7201), .Y(n7203) );
  OAI21XL U8814 ( .A0(n3421), .A1(n8275), .B0(n7204), .Y(n7206) );
  OAI21XL U8815 ( .A0(n7956), .A1(n8282), .B0(n7207), .Y(n7209) );
  OAI21XL U8816 ( .A0(n3359), .A1(n8387), .B0(n7210), .Y(n7212) );
  OAI21XL U8817 ( .A0(n7963), .A1(n8289), .B0(n7213), .Y(n7215) );
  OAI21XL U8818 ( .A0(n7068), .A1(n8289), .B0(n7216), .Y(n7218) );
  OAI21XL U8819 ( .A0(n7963), .A1(n8387), .B0(n7219), .Y(n7221) );
  OAI21XL U8820 ( .A0(n7068), .A1(n8125), .B0(n7222), .Y(n7224) );
  OAI21XL U8821 ( .A0(n7963), .A1(n8125), .B0(n7225), .Y(n7227) );
  OAI21XL U8822 ( .A0(n7956), .A1(n8387), .B0(n7228), .Y(n7230) );
  OAI21XL U8823 ( .A0(n3359), .A1(n8425), .B0(n7231), .Y(n7233) );
  OAI21XL U8824 ( .A0(n3421), .A1(n8387), .B0(n7234), .Y(n7236) );
  OAI21XL U8825 ( .A0(n3374), .A1(n8289), .B0(n7237), .Y(n7239) );
  OAI21XL U8826 ( .A0(n3391), .A1(n8289), .B0(n7240), .Y(n7242) );
  OAI21XL U8827 ( .A0(n3391), .A1(n8381), .B0(n7243), .Y(n7245) );
  OAI21XL U8828 ( .A0(n7068), .A1(n8310), .B0(n7246), .Y(n7248) );
  OAI21XL U8829 ( .A0(n7956), .A1(n8130), .B0(n7249), .Y(n7251) );
  OAI21XL U8830 ( .A0(n7068), .A1(n8317), .B0(n7252), .Y(n7254) );
  OAI21XL U8831 ( .A0(n3391), .A1(n8136), .B0(n7255), .Y(n7257) );
  OAI21XL U8832 ( .A0(n3359), .A1(n8349), .B0(n7258), .Y(n7260) );
  OAI21XL U8833 ( .A0(n7956), .A1(n3405), .B0(n7262), .Y(n7264) );
  OAI21XL U8834 ( .A0(n7963), .A1(n8349), .B0(n7265), .Y(n7267) );
  OAI21XL U8835 ( .A0(n3391), .A1(n7907), .B0(n7268), .Y(n7270) );
  OAI21XL U8836 ( .A0(n3374), .A1(n7907), .B0(n7271), .Y(n7273) );
  OAI21XL U8837 ( .A0(n3374), .A1(n3397), .B0(n7274), .Y(n7276) );
  OAI21XL U8838 ( .A0(n3391), .A1(n3397), .B0(n7277), .Y(n7279) );
  OAI21XL U8839 ( .A0(n3374), .A1(n8454), .B0(n7280), .Y(n7282) );
  OAI21XL U8840 ( .A0(n3391), .A1(n8454), .B0(n7283), .Y(n7285) );
  OAI21XL U8841 ( .A0(n3374), .A1(n8387), .B0(n7286), .Y(n7288) );
  OAI21XL U8842 ( .A0(n3359), .A1(n7918), .B0(n7289), .Y(n7291) );
  OAI21XL U8843 ( .A0(n3391), .A1(n8387), .B0(n7292), .Y(n7294) );
  OAI21XL U8844 ( .A0(n7963), .A1(n7918), .B0(n7295), .Y(n7297) );
  OAI21XL U8845 ( .A0(n3421), .A1(n7907), .B0(n7299), .Y(n7301) );
  OAI21XL U8846 ( .A0(n7956), .A1(n7907), .B0(n7302), .Y(n7305) );
  OAI21XL U8847 ( .A0(n7307), .A1(n7306), .B0(n7303), .Y(n7310) );
  OAI21XL U8848 ( .A0(n3391), .A1(n3405), .B0(n7308), .Y(n7309) );
  OAI21XL U8849 ( .A0(n8035), .A1(n8282), .B0(n7313), .Y(n7315) );
  OAI21XL U8850 ( .A0(n3419), .A1(n7317), .B0(n7316), .Y(n7319) );
  OAI21XL U8851 ( .A0(n3385), .A1(n8136), .B0(n7320), .Y(n7322) );
  OAI21XL U8852 ( .A0(n8055), .A1(n8136), .B0(n7323), .Y(n7325) );
  OAI21XL U8853 ( .A0(n3370), .A1(n3397), .B0(n7327), .Y(n7329) );
  OAI21XL U8854 ( .A0(n3370), .A1(n8351), .B0(n7330), .Y(n7332) );
  OAI21XL U8855 ( .A0(n8055), .A1(n8153), .B0(n7333), .Y(n7335) );
  OAI21XL U8856 ( .A0(n3419), .A1(n8171), .B0(n7336), .Y(n7338) );
  OAI21XL U8857 ( .A0(n3370), .A1(n8165), .B0(n7339), .Y(n7341) );
  OAI21XL U8858 ( .A0(n3385), .A1(n8393), .B0(n7342), .Y(n7344) );
  OAI21XL U8859 ( .A0(n3419), .A1(n8329), .B0(n7345), .Y(n7347) );
  OAI21XL U8860 ( .A0(n3370), .A1(n8329), .B0(n7348), .Y(n7351) );
  OAI21XL U8861 ( .A0(n3370), .A1(n8159), .B0(n7353), .Y(n7355) );
  OAI21XL U8862 ( .A0(n3419), .A1(n8165), .B0(n7356), .Y(n7358) );
  OAI21XL U8863 ( .A0(n3419), .A1(n8159), .B0(n7359), .Y(n7361) );
  OAI21XL U8864 ( .A0(n3370), .A1(n8171), .B0(n7362), .Y(n7364) );
  OAI21XL U8865 ( .A0(n8055), .A1(n8406), .B0(n7365), .Y(n7367) );
  OAI21XL U8866 ( .A0(n3385), .A1(n8406), .B0(n7368), .Y(n7370) );
  OAI21XL U8867 ( .A0(n8323), .A1(n8035), .B0(n7371), .Y(n7373) );
  OAI21XL U8868 ( .A0(n8055), .A1(n8304), .B0(n7374), .Y(n7376) );
  OAI21XL U8869 ( .A0(n8035), .A1(n8425), .B0(n7378), .Y(n7380) );
  OAI21XL U8870 ( .A0(n3385), .A1(n8267), .B0(n7381), .Y(n7383) );
  OAI21XL U8871 ( .A0(n3370), .A1(n8217), .B0(n7384), .Y(n7386) );
  OAI21XL U8872 ( .A0(n3419), .A1(n3405), .B0(n7387), .Y(n7389) );
  OAI21XL U8873 ( .A0(n3370), .A1(n8202), .B0(n7390), .Y(n7392) );
  OAI21XL U8874 ( .A0(n8035), .A1(n7975), .B0(n7393), .Y(n7395) );
  OAI21XL U8875 ( .A0(n3419), .A1(n8202), .B0(n7396), .Y(n7398) );
  OAI21XL U8876 ( .A0(n8111), .A1(n7975), .B0(n7399), .Y(n7401) );
  OAI21XL U8877 ( .A0(n3385), .A1(n8209), .B0(n7402), .Y(n7404) );
  OAI21XL U8878 ( .A0(n7445), .A1(n8304), .B0(n7405), .Y(n7407) );
  OAI21XL U8879 ( .A0(n3385), .A1(n3397), .B0(n7408), .Y(n7410) );
  OAI21XL U8880 ( .A0(n3370), .A1(n8381), .B0(n7411), .Y(n7413) );
  OAI21XL U8881 ( .A0(n8055), .A1(n8159), .B0(n7414), .Y(n7416) );
  OAI21XL U8882 ( .A0(n8055), .A1(n3397), .B0(n7417), .Y(n7419) );
  OAI21XL U8883 ( .A0(n7507), .A1(n8432), .B0(n7420), .Y(n7422) );
  OAI21XL U8884 ( .A0(n8055), .A1(n8351), .B0(n7423), .Y(n7425) );
  OAI21XL U8885 ( .A0(n3385), .A1(n8351), .B0(n7426), .Y(n7428) );
  OAI21XL U8886 ( .A0(n8035), .A1(n7684), .B0(n7429), .Y(n7431) );
  OAI21XL U8887 ( .A0(n7445), .A1(n8425), .B0(n7432), .Y(n7434) );
  OAI21XL U8888 ( .A0(n3385), .A1(n7995), .B0(n7435), .Y(n7437) );
  OAI21XL U8889 ( .A0(n8055), .A1(n7995), .B0(n7438), .Y(n7440) );
  OAI21XL U8890 ( .A0(n3370), .A1(n7455), .B0(n7441), .Y(n7443) );
  OAI21XL U8891 ( .A0(n7445), .A1(n8275), .B0(n7444), .Y(n7447) );
  OAI21XL U8892 ( .A0(n8055), .A1(n8275), .B0(n7448), .Y(n7450) );
  OAI21XL U8893 ( .A0(n3370), .A1(n8267), .B0(n7451), .Y(n7453) );
  OAI21XL U8894 ( .A0(n3419), .A1(n7455), .B0(n7454), .Y(n7457) );
  OAI21XL U8895 ( .A0(n3419), .A1(n8387), .B0(n7458), .Y(n7460) );
  OAI21XL U8896 ( .A0(n3419), .A1(n8289), .B0(n7461), .Y(n7463) );
  OAI21XL U8897 ( .A0(n3370), .A1(n8387), .B0(n7464), .Y(n7466) );
  OAI21XL U8898 ( .A0(n3370), .A1(n8289), .B0(n7467), .Y(n7469) );
  OAI21XL U8899 ( .A0(n3419), .A1(n8125), .B0(n7470), .Y(n7472) );
  OAI21XL U8900 ( .A0(n3370), .A1(n8125), .B0(n7473), .Y(n7475) );
  OAI21XL U8901 ( .A0(n3385), .A1(n8387), .B0(n7476), .Y(n7478) );
  OAI21XL U8902 ( .A0(n8055), .A1(n8387), .B0(n7479), .Y(n7481) );
  OAI21XL U8903 ( .A0(n8111), .A1(n8289), .B0(n7482), .Y(n7485) );
  OAI21XL U8904 ( .A0(n8035), .A1(n8381), .B0(n7488), .Y(n7490) );
  OAI21XL U8905 ( .A0(n8111), .A1(n8381), .B0(n7491), .Y(n7493) );
  OAI21XL U8906 ( .A0(n3419), .A1(n8317), .B0(n7494), .Y(n7496) );
  OAI21XL U8907 ( .A0(n3419), .A1(n8310), .B0(n7497), .Y(n7499) );
  OAI21XL U8908 ( .A0(n3370), .A1(n8310), .B0(n7500), .Y(n7502) );
  OAI21XL U8909 ( .A0(n3370), .A1(n8282), .B0(n7503), .Y(n7505) );
  OAI21XL U8910 ( .A0(n3419), .A1(n8282), .B0(n7506), .Y(n7509) );
  OAI21XL U8911 ( .A0(n3419), .A1(n8070), .B0(n7510), .Y(n7512) );
  OAI21XL U8912 ( .A0(n8035), .A1(n8125), .B0(n7514), .Y(n7516) );
  OAI21XL U8913 ( .A0(n3419), .A1(n8370), .B0(n7518), .Y(n7520) );
  OAI21XL U8914 ( .A0(n8055), .A1(n8171), .B0(n7521), .Y(n7523) );
  OAI21XL U8915 ( .A0(n8111), .A1(n8351), .B0(n7524), .Y(n7526) );
  OAI21XL U8916 ( .A0(n3385), .A1(n7975), .B0(n7527), .Y(n7529) );
  OAI21XL U8917 ( .A0(n8111), .A1(n3397), .B0(n7530), .Y(n7532) );
  OAI21XL U8918 ( .A0(n8035), .A1(n3397), .B0(n7533), .Y(n7535) );
  OAI21XL U8919 ( .A0(n8055), .A1(n7620), .B0(n7536), .Y(n7538) );
  OAI21XL U8920 ( .A0(n3385), .A1(n7620), .B0(n7539), .Y(n7541) );
  OAI21XL U8921 ( .A0(n8111), .A1(n8387), .B0(n7542), .Y(n7544) );
  OAI21XL U8922 ( .A0(n3419), .A1(n7918), .B0(n7545), .Y(n7547) );
  OAI21XL U8923 ( .A0(n3370), .A1(n7918), .B0(n7548), .Y(n7550) );
  OAI21XL U8924 ( .A0(n8035), .A1(n8387), .B0(n7551), .Y(n7553) );
  OAI21XL U8925 ( .A0(n3385), .A1(n7907), .B0(n7554), .Y(n7556) );
  OAI21XL U8926 ( .A0(n3370), .A1(n7925), .B0(n7557), .Y(n7559) );
  OAI21XL U8927 ( .A0(n7578), .A1(n7560), .B0(n6959), .Y(n7563) );
  OAI21XL U8928 ( .A0(n3393), .A1(n8101), .B0(n7561), .Y(n7562) );
  OAI21XL U8929 ( .A0(n3394), .A1(n3397), .B0(n6959), .Y(n7568) );
  OAI21XL U8930 ( .A0(n7578), .A1(n7566), .B0(n7565), .Y(n7567) );
  OAI21XL U8931 ( .A0(n7570), .A1(n8406), .B0(n6959), .Y(n7574) );
  OAI21XL U8932 ( .A0(n7578), .A1(n7572), .B0(n7571), .Y(n7573) );
  OAI21XL U8933 ( .A0(n3393), .A1(n8130), .B0(n6959), .Y(n7580) );
  OAI21XL U8934 ( .A0(n7578), .A1(n7577), .B0(n7576), .Y(n7579) );
  OAI21XL U8935 ( .A0(n7740), .A1(n3399), .B0(n7586), .Y(n7588) );
  OAI21XL U8936 ( .A0(n3396), .A1(n8406), .B0(n7589), .Y(n7591) );
  OAI21XL U8937 ( .A0(n3396), .A1(n8393), .B0(n7592), .Y(n7594) );
  OAI21XL U8938 ( .A0(n3392), .A1(n8446), .B0(n7595), .Y(n7597) );
  OAI21XL U8939 ( .A0(n3396), .A1(n7995), .B0(n7598), .Y(n7600) );
  OAI21XL U8940 ( .A0(n8432), .A1(n3392), .B0(n7601), .Y(n7603) );
  OAI21XL U8941 ( .A0(n7740), .A1(n8387), .B0(n7604), .Y(n7606) );
  OAI21XL U8942 ( .A0(n3392), .A1(n8419), .B0(n7607), .Y(n7609) );
  OAI21XL U8943 ( .A0(n3396), .A1(n3399), .B0(n7610), .Y(n7612) );
  OAI21XL U8944 ( .A0(n7740), .A1(n8425), .B0(n7613), .Y(n7615) );
  OAI21XL U8945 ( .A0(n3396), .A1(n8323), .B0(n7616), .Y(n7618) );
  OAI21XL U8946 ( .A0(n5812), .A1(n7620), .B0(n7619), .Y(n7622) );
  OAI21XL U8947 ( .A0(n3392), .A1(n8282), .B0(n7623), .Y(n7625) );
  OAI21XL U8948 ( .A0(n3392), .A1(n8130), .B0(n7626), .Y(n7628) );
  OAI21XL U8949 ( .A0(n3396), .A1(n8153), .B0(n7629), .Y(n7631) );
  OAI21XL U8950 ( .A0(n7740), .A1(n3397), .B0(n7632), .Y(n7634) );
  OAI21XL U8951 ( .A0(n7740), .A1(n8351), .B0(n7635), .Y(n7637) );
  OAI21XL U8952 ( .A0(n3396), .A1(n8136), .B0(n7638), .Y(n7640) );
  OAI21XL U8953 ( .A0(n7740), .A1(n7907), .B0(n7641), .Y(n7643) );
  OAI21XL U8954 ( .A0(n7740), .A1(n8159), .B0(n7644), .Y(n7646) );
  OAI21XL U8955 ( .A0(n3392), .A1(n8209), .B0(n7647), .Y(n7649) );
  OAI21XL U8956 ( .A0(n3392), .A1(n8310), .B0(n7650), .Y(n7652) );
  OAI21XL U8957 ( .A0(n3396), .A1(n8209), .B0(n7653), .Y(n7655) );
  OAI21XL U8958 ( .A0(n3396), .A1(n8370), .B0(n7656), .Y(n7658) );
  OAI21XL U8959 ( .A0(n3392), .A1(n7975), .B0(n7659), .Y(n7661) );
  OAI21XL U8960 ( .A0(n3392), .A1(n8393), .B0(n7662), .Y(n7664) );
  OAI21XL U8961 ( .A0(n7740), .A1(n8381), .B0(n7665), .Y(n7667) );
  OAI21XL U8962 ( .A0(n7740), .A1(n8432), .B0(n7668), .Y(n7670) );
  OAI21XL U8963 ( .A0(n7740), .A1(n8076), .B0(n7671), .Y(n7673) );
  OAI21XL U8964 ( .A0(n7740), .A1(n3405), .B0(n7674), .Y(n7676) );
  OAI21XL U8965 ( .A0(n5812), .A1(n3397), .B0(n7677), .Y(n7679) );
  OAI21XL U8966 ( .A0(n3396), .A1(n8351), .B0(n7680), .Y(n7682) );
  OAI21XL U8967 ( .A0(n3392), .A1(n7684), .B0(n7683), .Y(n7686) );
  OAI21XL U8968 ( .A0(n5812), .A1(n8275), .B0(n7687), .Y(n7689) );
  OAI21XL U8969 ( .A0(n3396), .A1(n8282), .B0(n7691), .Y(n7693) );
  OAI21XL U8970 ( .A0(n7740), .A1(n8289), .B0(n7694), .Y(n7696) );
  OAI21XL U8971 ( .A0(n7740), .A1(n8125), .B0(n7697), .Y(n7700) );
  OAI21XL U8972 ( .A0(n7740), .A1(n8177), .B0(n7702), .Y(n7704) );
  OAI21XL U8973 ( .A0(n3392), .A1(n8381), .B0(n7705), .Y(n7707) );
  OAI21XL U8974 ( .A0(n7740), .A1(n8310), .B0(n7708), .Y(n7710) );
  OAI21XL U8975 ( .A0(n3396), .A1(n8217), .B0(n7711), .Y(n7713) );
  OAI21XL U8976 ( .A0(n3396), .A1(n8130), .B0(n7714), .Y(n7716) );
  OAI21XL U8977 ( .A0(n7740), .A1(n8282), .B0(n7717), .Y(n7719) );
  OAI21XL U8978 ( .A0(n3396), .A1(n8381), .B0(n7720), .Y(n7722) );
  OAI21XL U8979 ( .A0(n7740), .A1(n8370), .B0(n7724), .Y(n7726) );
  OAI21XL U8980 ( .A0(n7740), .A1(n8349), .B0(n7727), .Y(n7729) );
  OAI21XL U8981 ( .A0(n3396), .A1(n7975), .B0(n7730), .Y(n7732) );
  OAI21XL U8982 ( .A0(n3392), .A1(n3397), .B0(n7733), .Y(n7735) );
  OAI21XL U8983 ( .A0(n3392), .A1(n8387), .B0(n7736), .Y(n7738) );
  OAI21XL U8984 ( .A0(n7740), .A1(n7918), .B0(n7739), .Y(n7742) );
  OAI21XL U8985 ( .A0(n5812), .A1(n7907), .B0(n7743), .Y(n7745) );
  OAI21XL U8986 ( .A0(n3372), .A1(n7995), .B0(n7751), .Y(n7753) );
  OAI21XL U8987 ( .A0(n7773), .A1(n8370), .B0(n7755), .Y(n7757) );
  OAI21XL U8988 ( .A0(n7895), .A1(n8406), .B0(n7758), .Y(n7760) );
  OAI21XL U8989 ( .A0(n7773), .A1(n8446), .B0(n7762), .Y(n7764) );
  OAI21XL U8990 ( .A0(n7895), .A1(n7995), .B0(n7765), .Y(n7768) );
  OAI21XL U8991 ( .A0(n3372), .A1(n8387), .B0(n7770), .Y(n7772) );
  OAI21XL U8992 ( .A0(n7773), .A1(n8419), .B0(n7774), .Y(n7776) );
  OAI21XL U8993 ( .A0(n3372), .A1(n8393), .B0(n7777), .Y(n7779) );
  OAI21XL U8994 ( .A0(n7895), .A1(n8412), .B0(n7780), .Y(n7782) );
  OAI21XL U8995 ( .A0(n7773), .A1(n8412), .B0(n7783), .Y(n7785) );
  OAI21XL U8996 ( .A0(n7895), .A1(n8323), .B0(n7786), .Y(n7788) );
  OAI21XL U8997 ( .A0(n7773), .A1(n8454), .B0(n7789), .Y(n7791) );
  OAI21XL U8998 ( .A0(n7773), .A1(n8130), .B0(n7792), .Y(n7794) );
  OAI21XL U8999 ( .A0(n3372), .A1(n3397), .B0(n7796), .Y(n7798) );
  OAI21XL U9000 ( .A0(n3372), .A1(n8351), .B0(n7799), .Y(n7801) );
  OAI21XL U9001 ( .A0(n7895), .A1(n8136), .B0(n7802), .Y(n7804) );
  OAI21XL U9002 ( .A0(n7895), .A1(n8153), .B0(n7805), .Y(n7807) );
  OAI21XL U9003 ( .A0(n7895), .A1(n8393), .B0(n7808), .Y(n7810) );
  OAI21XL U9004 ( .A0(n7895), .A1(n8177), .B0(n7811), .Y(n7813) );
  OAI21XL U9005 ( .A0(n3372), .A1(n8171), .B0(n7814), .Y(n7816) );
  OAI21XL U9006 ( .A0(n3372), .A1(n8165), .B0(n7817), .Y(n7819) );
  OAI21XL U9007 ( .A0(n8323), .A1(n7773), .B0(n7820), .Y(n7822) );
  OAI21XL U9008 ( .A0(n7773), .A1(n8393), .B0(n7823), .Y(n7825) );
  OAI21XL U9009 ( .A0(n7773), .A1(n7975), .B0(n7827), .Y(n7829) );
  OAI21XL U9010 ( .A0(n3372), .A1(n8217), .B0(n7830), .Y(n7832) );
  OAI21XL U9011 ( .A0(n7895), .A1(n8304), .B0(n7833), .Y(n7835) );
  OAI21XL U9012 ( .A0(n7895), .A1(n8209), .B0(n7836), .Y(n7838) );
  OAI21XL U9013 ( .A0(n7895), .A1(n3397), .B0(n7839), .Y(n7841) );
  OAI21XL U9014 ( .A0(n3372), .A1(n8076), .B0(n7842), .Y(n7844) );
  OAI21XL U9015 ( .A0(n3372), .A1(n3405), .B0(n7845), .Y(n7847) );
  OAI21XL U9016 ( .A0(n3372), .A1(n8446), .B0(n7848), .Y(n7850) );
  OAI21XL U9017 ( .A0(n3372), .A1(n8381), .B0(n7851), .Y(n7853) );
  OAI21XL U9018 ( .A0(n7895), .A1(n8351), .B0(n7854), .Y(n7856) );
  OAI21XL U9019 ( .A0(n7895), .A1(n8425), .B0(n7857), .Y(n7859) );
  OAI21XL U9020 ( .A0(n7895), .A1(n8275), .B0(n7860), .Y(n7862) );
  OAI21XL U9021 ( .A0(n7773), .A1(n7864), .B0(n7863), .Y(n7866) );
  OAI21XL U9022 ( .A0(n3372), .A1(n8289), .B0(n7867), .Y(n7869) );
  OAI21XL U9023 ( .A0(n7895), .A1(n8387), .B0(n7870), .Y(n7872) );
  OAI21XL U9024 ( .A0(n7773), .A1(n8381), .B0(n7873), .Y(n7876) );
  OAI21XL U9025 ( .A0(n7773), .A1(n7878), .B0(n7877), .Y(n7880) );
  OAI21XL U9026 ( .A0(n3372), .A1(n8310), .B0(n7881), .Y(n7883) );
  OAI21XL U9027 ( .A0(n3372), .A1(n8323), .B0(n7884), .Y(n7886) );
  OAI21XL U9028 ( .A0(n3372), .A1(n8282), .B0(n7889), .Y(n7892) );
  OAI21XL U9029 ( .A0(n7895), .A1(n8381), .B0(n7894), .Y(n7897) );
  OAI21XL U9030 ( .A0(n3372), .A1(n8349), .B0(n7899), .Y(n7901) );
  OAI21XL U9031 ( .A0(n3372), .A1(n8370), .B0(n7903), .Y(n7905) );
  OAI21XL U9032 ( .A0(n7773), .A1(n7907), .B0(n7906), .Y(n7909) );
  OAI21XL U9033 ( .A0(n7773), .A1(n3397), .B0(n7911), .Y(n7913) );
  OAI21XL U9034 ( .A0(n7773), .A1(n8387), .B0(n7914), .Y(n7916) );
  OAI21XL U9035 ( .A0(n3372), .A1(n7918), .B0(n7917), .Y(n7921) );
  OAI21XL U9036 ( .A0(n3372), .A1(n7925), .B0(n7924), .Y(n7928) );
  OAI21XL U9037 ( .A0(n7956), .A1(n8419), .B0(n7943), .Y(n7945) );
  OAI21XL U9038 ( .A0(n3391), .A1(n8446), .B0(n7946), .Y(n7948) );
  OAI21XL U9039 ( .A0(n7956), .A1(n8432), .B0(n7949), .Y(n7951) );
  OAI21XL U9040 ( .A0(n3391), .A1(n8419), .B0(n7952), .Y(n7954) );
  OAI21XL U9041 ( .A0(n7956), .A1(n3399), .B0(n7955), .Y(n7958) );
  OAI21XL U9042 ( .A0(n3391), .A1(n8059), .B0(n7959), .Y(n7961) );
  OAI21XL U9043 ( .A0(n7963), .A1(n8425), .B0(n7962), .Y(n7965) );
  OAI21XL U9044 ( .A0(n3391), .A1(n8440), .B0(n7966), .Y(n7968) );
  OAI21XL U9045 ( .A0(n3391), .A1(n8412), .B0(n7969), .Y(n7971) );
  OAI21XL U9046 ( .A0(n3374), .A1(n8446), .B0(n7988), .Y(n7990) );
  OAI21XL U9047 ( .A0(n3374), .A1(n8419), .B0(n7991), .Y(n7993) );
  OAI21XL U9048 ( .A0(n3359), .A1(n7995), .B0(n7994), .Y(n7997) );
  OAI21XL U9049 ( .A0(n3421), .A1(n3399), .B0(n7998), .Y(n8000) );
  OAI21XL U9050 ( .A0(n3421), .A1(n8412), .B0(n8001), .Y(n8003) );
  OAI21XL U9051 ( .A0(n3374), .A1(n8370), .B0(n8004), .Y(n8006) );
  OAI21XL U9052 ( .A0(n8432), .A1(n3374), .B0(n8007), .Y(n8009) );
  OAI21XL U9053 ( .A0(n3421), .A1(n8323), .B0(n8010), .Y(n8012) );
  OAI21XL U9054 ( .A0(n3421), .A1(n8446), .B0(n8013), .Y(n8016) );
  OAI21XL U9055 ( .A0(n3374), .A1(n3399), .B0(n8017), .Y(n8020) );
  OAI21XL U9056 ( .A0(n8055), .A1(n8419), .B0(n8039), .Y(n8041) );
  OAI21XL U9057 ( .A0(n8055), .A1(n8059), .B0(n8042), .Y(n8044) );
  OAI21XL U9058 ( .A0(n8055), .A1(n8432), .B0(n8045), .Y(n8047) );
  OAI21XL U9059 ( .A0(n8035), .A1(n8446), .B0(n8048), .Y(n8050) );
  OAI21XL U9060 ( .A0(n8035), .A1(n8419), .B0(n8051), .Y(n8053) );
  OAI21XL U9061 ( .A0(n8055), .A1(n3399), .B0(n8054), .Y(n8057) );
  OAI21XL U9062 ( .A0(n8035), .A1(n8059), .B0(n8058), .Y(n8061) );
  OAI21XL U9063 ( .A0(n3370), .A1(n8425), .B0(n8062), .Y(n8064) );
  OAI21XL U9064 ( .A0(n3370), .A1(n8419), .B0(n8065), .Y(n8067) );
  OAI21XL U9065 ( .A0(n3385), .A1(n8432), .B0(n8085), .Y(n8088) );
  OAI21XL U9066 ( .A0(n3385), .A1(n3399), .B0(n8090), .Y(n8093) );
  OAI21XL U9067 ( .A0(n7507), .A1(n3399), .B0(n8095), .Y(n8098) );
  OAI21XL U9068 ( .A0(n3419), .A1(n8101), .B0(n8100), .Y(n8103) );
  OAI21XL U9069 ( .A0(n8111), .A1(n8419), .B0(n8104), .Y(n8106) );
  OAI21XL U9070 ( .A0(n8111), .A1(n8446), .B0(n8107), .Y(n8109) );
  OAI21XL U9071 ( .A0(n8432), .A1(n8111), .B0(n8110), .Y(n8113) );
  OAI21XL U9072 ( .A0(n3419), .A1(n8425), .B0(n8115), .Y(n8117) );
  OAI21XL U9073 ( .A0(n3385), .A1(n8323), .B0(n8118), .Y(n8120) );
  OAI21XL U9074 ( .A0(n3385), .A1(n8446), .B0(n8121), .Y(n8123) );
  OAI21XL U9075 ( .A0(n8447), .A1(n8125), .B0(n8124), .Y(n8127) );
  OAI21XL U9076 ( .A0(n6407), .A1(n8130), .B0(n8129), .Y(n8133) );
  OAI21XL U9077 ( .A0(n8447), .A1(n8136), .B0(n8135), .Y(n8139) );
  OAI21XL U9078 ( .A0(n3386), .A1(n8351), .B0(n8142), .Y(n8145) );
  OAI21XL U9079 ( .A0(n3386), .A1(n3397), .B0(n8147), .Y(n8150) );
  OAI21XL U9080 ( .A0(n8447), .A1(n8153), .B0(n8152), .Y(n8156) );
  OAI21XL U9081 ( .A0(n3386), .A1(n8159), .B0(n8158), .Y(n8162) );
  OAI21XL U9082 ( .A0(n8268), .A1(n8165), .B0(n8164), .Y(n8168) );
  OAI21XL U9083 ( .A0(n3386), .A1(n8171), .B0(n8170), .Y(n8174) );
  OAI21XL U9084 ( .A0(n8447), .A1(n8177), .B0(n8176), .Y(n8180) );
  OAI21XL U9085 ( .A0(n8268), .A1(n8184), .B0(n8183), .Y(n8187) );
  OAI21XL U9086 ( .A0(n8447), .A1(n8289), .B0(n8189), .Y(n8192) );
  OAI21XL U9087 ( .A0(n6407), .A1(n8425), .B0(n8194), .Y(n8197) );
  OAI21XL U9088 ( .A0(n3386), .A1(n8202), .B0(n8201), .Y(n8205) );
  OAI21XL U9089 ( .A0(n6407), .A1(n8209), .B0(n8208), .Y(n8212) );
  OAI21XL U9090 ( .A0(n3386), .A1(n8217), .B0(n8216), .Y(n8220) );
  OAI21XL U9091 ( .A0(n8268), .A1(n8381), .B0(n8223), .Y(n8226) );
  OAI21XL U9092 ( .A0(n6407), .A1(n8267), .B0(n8229), .Y(n8232) );
  OAI21XL U9093 ( .A0(n8447), .A1(n3397), .B0(n8234), .Y(n8237) );
  OAI21XL U9094 ( .A0(n8447), .A1(n8310), .B0(n8239), .Y(n8242) );
  OAI21XL U9095 ( .A0(n3386), .A1(n8432), .B0(n8244), .Y(n8247) );
  OAI21XL U9096 ( .A0(n3386), .A1(n8446), .B0(n8249), .Y(n8252) );
  OAI21XL U9097 ( .A0(n8447), .A1(n8351), .B0(n8254), .Y(n8257) );
  OAI21XL U9098 ( .A0(n3386), .A1(n8275), .B0(n8261), .Y(n8264) );
  OAI21XL U9099 ( .A0(n8268), .A1(n8267), .B0(n8266), .Y(n8271) );
  OAI21XL U9100 ( .A0(n8447), .A1(n8275), .B0(n8274), .Y(n8278) );
  OAI21XL U9101 ( .A0(n8447), .A1(n8282), .B0(n8281), .Y(n8285) );
  OAI21XL U9102 ( .A0(n3386), .A1(n8289), .B0(n8288), .Y(n8292) );
  OAI21XL U9103 ( .A0(n3386), .A1(n8412), .B0(n8296), .Y(n8299) );
  OAI21XL U9104 ( .A0(n6407), .A1(n8304), .B0(n8303), .Y(n8307) );
  OAI21XL U9105 ( .A0(n3386), .A1(n8310), .B0(n8309), .Y(n8313) );
  OAI21XL U9106 ( .A0(n3386), .A1(n8317), .B0(n8316), .Y(n8320) );
  OAI21XL U9107 ( .A0(n3386), .A1(n8323), .B0(n8322), .Y(n8326) );
  OAI21XL U9108 ( .A0(n8447), .A1(n8329), .B0(n8328), .Y(n8332) );
  OAI21XL U9109 ( .A0(n8447), .A1(n8381), .B0(n8335), .Y(n8338) );
  OAI21XL U9110 ( .A0(n3386), .A1(n8370), .B0(n8344), .Y(n8347) );
  OAI21XL U9111 ( .A0(n6407), .A1(n8351), .B0(n8350), .Y(n8354) );
  OAI21XL U9112 ( .A0(n6407), .A1(n3397), .B0(n8357), .Y(n8360) );
  OAI21XL U9113 ( .A0(n6407), .A1(n8387), .B0(n8363), .Y(n8366) );
  OAI21XL U9114 ( .A0(n3386), .A1(n8387), .B0(n8386), .Y(n8390) );
  OAI21XL U9115 ( .A0(n8447), .A1(n8393), .B0(n8392), .Y(n8396) );
  OAI21XL U9116 ( .A0(n6407), .A1(n8446), .B0(n8399), .Y(n8402) );
  OAI21XL U9117 ( .A0(n8447), .A1(n8406), .B0(n8405), .Y(n8409) );
  OAI21XL U9118 ( .A0(n8447), .A1(n8412), .B0(n8411), .Y(n8415) );
  OAI21XL U9119 ( .A0(n6407), .A1(n8419), .B0(n8418), .Y(n8422) );
  OAI21XL U9120 ( .A0(n3386), .A1(n8425), .B0(n8424), .Y(n8428) );
  OAI21XL U9121 ( .A0(n8432), .A1(n6407), .B0(n8431), .Y(n8435) );
  OAI21XL U9122 ( .A0(n6407), .A1(n8440), .B0(n8439), .Y(n8443) );
  OAI21XL U9123 ( .A0(n8447), .A1(n8446), .B0(n8445), .Y(n8450) );
  OAI21XL U9124 ( .A0(n6407), .A1(n8454), .B0(n8453), .Y(n8457) );
  ADDHXL U9125 ( .A(n8459), .B(n8458), .CO(DP_OP_2677J1_122_9848_n30), .S(
        n5259) );
  OAI21XL U9126 ( .A0(n8481), .A1(done), .B0(n8460), .Y(n3339) );
  OAI21XL U9127 ( .A0(n8534), .A1(n8463), .B0(n8462), .Y(n3343) );
  OAI21XL U9128 ( .A0(IROM_A[1]), .A1(n8465), .B0(n8464), .Y(n3338) );
  AOI22XL U9129 ( .A0(n8468), .A1(n8473), .B0(n8467), .B1(n8466), .Y(n8476) );
  OAI211XL U9130 ( .A0(n8472), .A1(n8471), .B0(n8470), .C0(n8469), .Y(n8485)
         );
  OAI21XL U9131 ( .A0(n8476), .A1(n8475), .B0(n8474), .Y(n3341) );
  AOI21XL U9132 ( .A0(n8480), .A1(in_done), .B0(n8566), .Y(n3340) );
  OAI21XL U9133 ( .A0(IROM_A[0]), .A1(n8478), .B0(n8477), .Y(n3333) );
  OAI21XL U9134 ( .A0(n8481), .A1(in_done), .B0(n8480), .Y(n3329) );
  AOI21XL U9135 ( .A0(n8483), .A1(op2[1]), .B0(n8482), .Y(n8484) );
  AOI21XL U9136 ( .A0(n8485), .A1(op2[1]), .B0(n8484), .Y(n3323) );
  OAI21XL U9137 ( .A0(IROM_A[3]), .A1(n8487), .B0(n8486), .Y(n3321) );
  AOI21XL U9138 ( .A0(IRAM_valid), .A1(n8489), .B0(n8488), .Y(n3320) );
  OAI21XL U9139 ( .A0(image_data[429]), .A1(n8498), .B0(n8497), .Y(n3237) );
  OAI21XL U9140 ( .A0(image_data[284]), .A1(n8507), .B0(n8506), .Y(n3092) );
  OAI21XL U9141 ( .A0(n8509), .A1(n8508), .B0(n3365), .Y(n8510) );
  OAI21XL U9142 ( .A0(n8515), .A1(n3417), .B0(n8514), .Y(n8516) );
  AOI21XL U9143 ( .A0(n3417), .A1(image_data[22]), .B0(n8516), .Y(n2830) );
endmodule

